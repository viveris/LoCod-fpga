-- 
-- Politecnico di Milano
-- Code created using PandA - Version: PandA 0.9.8 - Revision eda4c22d5adaec44fd8489ae49b854b244d2cf70-HEAD - Date 2023-03-02T09:23:24
-- bambu executed with: bambu --writer=H --generate-interface=MINIMAL --memory-allocation-policy=NO_BRAM --channels-type=MEM_ACC_11 --memory-ctrl-type=D21 --top-fname=acc_0 --top-rtldesign-name=acc_0 ../src/main.c 
-- 
-- Send any bug to: panda-info@polimi.it
-- ************************************************************************
-- The following text holds for all the components tagged with PANDA_LGPLv3.
-- They are all part of the BAMBU/PANDA IP LIBRARY.
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 3 of the License, or (at your option) any later version.
-- 
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
-- 
-- You should have received a copy of the GNU Lesser General Public
-- License along with the PandA framework; see the files COPYING.LIB
-- If not, see <http://www.gnu.org/licenses/>.
-- ************************************************************************


library IEEE;
use IEEE.numeric_std.all;

package panda_pkg is
   function resize_signed(input : signed; size : integer) return signed;
end;

package body panda_pkg is
   function resize_signed(input : signed; size : integer) return signed is
   begin
     if (size > input'length) then
       return resize(input, size);
     else
       return input(size-1+input'right downto input'right);
     end if;
   end function;
end package body;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>, Christian Pilato <christian.pilato@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity constant_value is 
generic(
 BITSIZE_out1: integer;
 value: std_logic_vector);
port (
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end constant_value;

architecture constant_value_arch of constant_value is
  begin
   out1 <= value;
end constant_value_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity register_SE is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  wenable : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end register_SE;

architecture register_SE_arch of register_SE is
  
  signal reg_out1 : std_logic_vector(BITSIZE_out1-1 downto 0) := (others => '0');
  begin
    out1 <= reg_out1;
    process(clock)
    begin
      if(clock'event and clock = '1') then
        if(wenable = '1') then
          reg_out1 <= in1;
        end if;
      end if;
    end process;

end register_SE_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity register_STD is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  wenable : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end register_STD;

architecture register_STD_arch of register_STD is
  
  signal reg_out1 : std_logic_vector(BITSIZE_out1-1 downto 0) := (others => '0');
  begin
  out1 <= reg_out1;
  process(clock)
  begin
    if(clock'event and clock = '1') then
      reg_out1 <= in1;
    end if;
  end process;

end register_STD_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity UUdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end UUdata_converter_FU;

architecture UUdata_converter_FU_arch of UUdata_converter_FU is
  begin
  out1 <= std_logic_vector(resize(unsigned(in1), BITSIZE_out1));
end UUdata_converter_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2020-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity extract_bit_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out std_logic

);
end extract_bit_expr_FU;

architecture extract_bit_expr_FU_arch of extract_bit_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= shift_right(in1, to_integer(unsigned(in2)))(0);
    end process;

end extract_bit_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity IUdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end IUdata_converter_FU;

architecture IUdata_converter_FU_arch of IUdata_converter_FU is
  begin
    process(in1)
    begin
      if(BITSIZE_out1 <= BITSIZE_in1) then
        out1 <= unsigned(in1(BITSIZE_out1-1 downto 0));
      else
        out1 <= unsigned(resize(in1, BITSIZE_out1));
      end if;
    end process;
end IUdata_converter_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2016-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity lut_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  in2 : in std_logic;
  in3 : in std_logic;
  in4 : in std_logic;
  in5 : in std_logic;
  in6 : in std_logic;
  in7 : in std_logic;
  in8 : in std_logic;
  in9 : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end lut_expr_FU;

architecture lut_expr_FU_arch of lut_expr_FU is
    signal in0 : std_logic_vector(7 downto 0);
    signal shifted_s : unsigned(in1'range) := (others => '0');
  begin
    in0(0) <= in2;
    in0(1) <= in3;
    in0(2) <= in4;
    in0(3) <= in5;
    in0(4) <= in6;
    in0(5) <= in7;
    in0(6) <= in8;
    in0(7) <= in9;
    out1 <= std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (shifted_s(0) = '1') else (others => '0');
    process(in0, in1)
    begin
      shifted_s <= shift_right(unsigned(in1), to_integer(unsigned(in0)));
    end process;

end lut_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity UIdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end UIdata_converter_FU;

architecture UIdata_converter_FU_arch of UIdata_converter_FU is
  begin
    process(in1)
    begin
      if(BITSIZE_out1 > BITSIZE_in1) then
        out1 <= signed(resize(in1, BITSIZE_out1));
      else
        out1 <= signed(in1 (BITSIZE_out1-1 downto 0));
      end if;
    end process;
end UIdata_converter_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity IIdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end IIdata_converter_FU;

architecture IIdata_converter_FU_arch of IIdata_converter_FU is
  begin
    process(in1)
    begin
      if(BITSIZE_out1 > BITSIZE_in1) then
        out1 <= resize(in1, BITSIZE_out1);
      else
        out1 <= in1 (BITSIZE_out1-1 downto 0);
      end if;
    end process;
end IIdata_converter_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity multi_read_cond_FU is 
generic(
 BITSIZE_in1: integer;
 PORTSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end multi_read_cond_FU;

architecture multi_read_cond_FU_arch of multi_read_cond_FU is
  begin
    out1 <= in1;
end multi_read_cond_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2020-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_extract_bit_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out std_logic

);
end ui_extract_bit_expr_FU;

architecture ui_extract_bit_expr_FU_arch of ui_extract_bit_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= shift_right(unsigned(in1), to_integer(unsigned(in2)))(0);
    end process;

end ui_extract_bit_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bit_and_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end bit_and_expr_FU;

architecture bit_and_expr_FU_arch of bit_and_expr_FU is
  begin
  out1 <= resize_signed(in1, BITSIZE_out1) and resize_signed(in2, BITSIZE_out1);
end bit_and_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bit_ior_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end bit_ior_expr_FU;

architecture bit_ior_expr_FU_arch of bit_ior_expr_FU is
  begin
  out1 <= resize_signed(in1, BITSIZE_out1) or resize_signed(in2, BITSIZE_out1);
end bit_ior_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bit_not_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end bit_not_expr_FU;

architecture bit_not_expr_FU_arch of bit_not_expr_FU is
  begin
  out1 <= not resize_signed(in1, BITSIZE_out1);
end bit_not_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity eq_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end eq_expr_FU;

architecture eq_expr_FU_arch of eq_expr_FU is
  begin
    out1 <= std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (in1 = in2) else (others => '0');

end eq_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity minus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end minus_expr_FU;

architecture minus_expr_FU_arch of minus_expr_FU is
  begin
  out1 <= resize_signed(in1, BITSIZE_out1) - resize_signed(in2, BITSIZE_out1);
end minus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity mult_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PIPE_PARAMETER: integer);
port (
  -- IN
  clock : in std_logic;
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end mult_expr_FU;

architecture mult_expr_FU_arch of mult_expr_FU is
    signal in1_int : signed (BITSIZE_in1-1 downto 0);
    signal in2_int : signed (BITSIZE_in2-1 downto 0);
  begin
    cond: if(PIPE_PARAMETER=0) generate
      out1 <= signed(resize_signed(in1 * in2, BITSIZE_out1));
    end generate cond;
    cond1 : if(PIPE_PARAMETER=1) generate
      out1 <= resize_signed(in1_int * in2_int, BITSIZE_out1);
      process(clock)
      begin
        if clock'event and clock = '1' then
          in1_int <= resize(in1, BITSIZE_in1);
          in2_int <= resize(in2, BITSIZE_in2);
        end if;
      end process;
    end generate cond1;
    cond2 : if(PIPE_PARAMETER >1) generate
      type levels_of_registers is array (PIPE_PARAMETER-2 downto 0) of signed(BITSIZE_out1-1 downto 0);
      signal out1_int : levels_of_registers;
    begin
      process(clock)
      begin
        if clock'event and clock = '1' then
          in1_int <= in1;
          in2_int <= in2;
          out1_int(PIPE_PARAMETER-2) <= signed(resize_signed(signed(in1_int * in2_int), BITSIZE_out1));
          for i in 0 to PIPE_PARAMETER-3 loop
            out1_int (i) <= out1_int (i+1);
          end loop;
        end if;
      end process;
      out1 <= out1_int (0);
    end generate cond2;

end mult_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity negate_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end negate_expr_FU;

architecture negate_expr_FU_arch of negate_expr_FU is
  begin
    out1 <= -resize_signed(in1, BITSIZE_out1);

end negate_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity plus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end plus_expr_FU;

architecture plus_expr_FU_arch of plus_expr_FU is
    signal resized_in1 : signed (BITSIZE_out1-1 downto 0);
    signal resized_in2 : signed (BITSIZE_out1-1 downto 0);
    begin
      process(in1,in2,resized_in1,resized_in2)
      begin
        if(BITSIZE_out1 <= BITSIZE_in1) then
          resized_in1 <= in1(BITSIZE_out1-1 downto 0);
        else
          resized_in1 <= resize(in1, BITSIZE_out1);
        end if;
        if(BITSIZE_out1 < BITSIZE_in2) then
          resized_in2 <= in2(BITSIZE_out1-1 downto 0);
        else
          resized_in2 <= resize(in2, BITSIZE_out1);
        end if;
        out1 <= resized_in1 + resized_in2;
      end process;

end plus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_bit_and_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_bit_and_expr_FU;

architecture ui_bit_and_expr_FU_arch of ui_bit_and_expr_FU is
  begin
  out1 <= resize(in1, BITSIZE_out1) and resize(in2, BITSIZE_out1);
end ui_bit_and_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2016-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_bit_ior_concat_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_in3: integer;
 BITSIZE_out1: integer;
 OFFSET_PARAMETER: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  in3 : in unsigned (BITSIZE_in3-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_bit_ior_concat_expr_FU;

architecture ui_bit_ior_concat_expr_FU_arch of ui_bit_ior_concat_expr_FU is
  function integer_ternary_operator(cond : boolean; op1 : integer; op2 : integer) return integer is
    begin
      if cond then
        return op1;
      else
        return op2;
      end if;
  end integer_ternary_operator;
    constant nbit_out : integer := integer_ternary_operator(BITSIZE_out1 > OFFSET_PARAMETER, BITSIZE_out1, 1+OFFSET_PARAMETER);
    signal tmp_in1 : unsigned(nbit_out-1 downto 0);
    signal tmp_in2 : unsigned(nbit_out-1 downto 0);
    begin
      tmp_in1 <= resize(in1, nbit_out);
      tmp_in2 <= resize(in2, nbit_out);
      out1 <= resize(tmp_in1(nbit_out-1 downto OFFSET_PARAMETER) & tmp_in2(OFFSET_PARAMETER-1 downto 0), BITSIZE_out1);
      
end ui_bit_ior_concat_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_bit_ior_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_bit_ior_expr_FU;

architecture ui_bit_ior_expr_FU_arch of ui_bit_ior_expr_FU is
  begin
  out1 <= resize(in1, BITSIZE_out1) or resize(in2, BITSIZE_out1);
end ui_bit_ior_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_cond_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_in3: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  in3 : in unsigned (BITSIZE_in3-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_cond_expr_FU;

architecture ui_cond_expr_FU_arch of ui_cond_expr_FU is
  constant zeroes : std_logic_vector(in1'range) := (others => '0');
  begin
    out1 <= resize(in2, BITSIZE_out1) when (in1 /= zeroes) else resize(in3, BITSIZE_out1);

end ui_cond_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_eq_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end ui_eq_expr_FU;

architecture ui_eq_expr_FU_arch of ui_eq_expr_FU is
  begin
    out1 <= std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (in1 = in2) else (others => '0');

end ui_eq_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_lshift_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PRECISION: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_lshift_expr_FU;

architecture ui_lshift_expr_FU_arch of ui_lshift_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= shift_left(resize(in1, BITSIZE_out1), to_integer(unsigned(in2) rem PRECISION));
    end process;

end ui_lshift_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_mult_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PIPE_PARAMETER: integer);
port (
  -- IN
  clock : in std_logic;
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_mult_expr_FU;

architecture ui_mult_expr_FU_arch of ui_mult_expr_FU is
    signal in1_int : unsigned (BITSIZE_in1-1 downto 0);
    signal in2_int : unsigned (BITSIZE_in2-1 downto 0);
  begin
    cond: if(PIPE_PARAMETER=0) generate
      out1 <= resize(in1 * in2, BITSIZE_out1);
    end generate cond;
    cond1 : if(PIPE_PARAMETER=1) generate
      out1 <= resize(in1_int * in2_int, BITSIZE_out1);
      process(clock)
      begin
        if clock'event and clock = '1' then
          in1_int <= in1;
          in2_int <= in2;
        end if;
      end process;
    end generate cond1;
    cond2 : if(PIPE_PARAMETER >1) generate
      type levels_of_registers is array (PIPE_PARAMETER-1 downto 0) of unsigned (BITSIZE_out1-1 downto 0);
      signal out1_int : levels_of_registers;
    begin
      out1 <= out1_int (0);
      process(clock)
      begin
        if clock'event and clock = '1' then
          in1_int <= in1;
          in2_int <= in2;
          out1_int(PIPE_PARAMETER-2) <= resize(in1_int * in2_int, BITSIZE_out1);
          for i in 0 to PIPE_PARAMETER-3 loop
            out1_int (i) <= out1_int (i+1);
          end loop;
        end if;
      end process;
    end generate cond2;

end ui_mult_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_ne_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end ui_ne_expr_FU;

architecture ui_ne_expr_FU_arch of ui_ne_expr_FU is
  signal xs1 : unsigned(in1'range) := (others => 'X');
  signal xs2 : unsigned(in2'range) := (others => 'X');
  begin
    out1 <= (others => 'X') when (not((in1 >= in2) or (in1 <= in2))) else std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (in1 /= in2) else (others => '0');

end ui_ne_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_plus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_plus_expr_FU;

architecture ui_plus_expr_FU_arch of ui_plus_expr_FU is
    signal resized_in1 : unsigned(BITSIZE_out1-1 downto 0);
    signal resized_in2 : unsigned(BITSIZE_out1-1 downto 0);
    begin
      process(in1,in2,resized_in1,resized_in2)
      begin
        if(BITSIZE_out1 <= BITSIZE_in1) then
          resized_in1 <= in1(BITSIZE_out1-1 downto 0);
        else
          resized_in1 <= resize(in1, BITSIZE_out1);
        end if;
        if(BITSIZE_out1 < BITSIZE_in2) then
          resized_in2 <= in2(BITSIZE_out1-1 downto 0);
        else
          resized_in2 <= resize(in2, BITSIZE_out1);
        end if;
        out1 <= resized_in1 + resized_in2;
      end process;

end ui_plus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_pointer_plus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 LSB_PARAMETER: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_pointer_plus_expr_FU;

architecture ui_pointer_plus_expr_FU_arch of ui_pointer_plus_expr_FU is
  begin
    out1 <= resize(in1, BITSIZE_out1) + resize(in2, BITSIZE_out1);
end ui_pointer_plus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_rshift_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PRECISION: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_rshift_expr_FU;

architecture ui_rshift_expr_FU_arch of ui_rshift_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= resize(shift_right(in1, to_integer(unsigned(in2) rem PRECISION)), BITSIZE_out1);
    end process;

end ui_rshift_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_ternary_plus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_in3: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  in3 : in unsigned (BITSIZE_in3-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end ui_ternary_plus_expr_FU;

architecture ui_ternary_plus_expr_FU_arch of ui_ternary_plus_expr_FU is
  begin
  out1 <= resize(in1, BITSIZE_out1) + resize(in2, BITSIZE_out1) + resize(in3, BITSIZE_out1);
end ui_ternary_plus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2013-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bus_merger is 
generic(
 BITSIZE_in1: integer;
 PORTSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end bus_merger;

architecture bus_merger_arch of bus_merger is
  begin
  process(in1)
  variable temp_out1 : std_logic_vector(BITSIZE_out1-1 downto 0);
  begin
    temp_out1 := (others => '0');
    for I in 0 to PORTSIZE_in1-1 loop
      temp_out1 := temp_out1 or in1(((I+1)*BITSIZE_in1)-1 downto (I*BITSIZE_in1));
    end loop;  out1 <= temp_out1;
  end process;

end bus_merger_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ASSIGN_VECTOR_BOOL_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end ASSIGN_VECTOR_BOOL_FU;

architecture ASSIGN_VECTOR_BOOL_FU_arch of ASSIGN_VECTOR_BOOL_FU is
  begin
    out1 <= in1;
end ASSIGN_VECTOR_BOOL_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>, Christian Pilato <christian.pilato@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity MUX_GATE is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  sel : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end MUX_GATE;

architecture MUX_GATE_arch of MUX_GATE is
  begin
  out1 <= in1 when sel='1' else in2;
end MUX_GATE_arch;

-- Datapath RTL description for acc_0
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity datapath_acc_0 is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in_port_param : in std_logic_vector(31 downto 0) ;
  in_port_result : in std_logic_vector(31 downto 0) ;
  M_Rdata_ram : in std_logic_vector(31 downto 0) ;
  M_DataRdy : in std_logic;
  Min_oe_ram : in std_logic;
  Min_we_ram : in std_logic;
  Min_addr_ram : in std_logic_vector(31 downto 0) ;
  Min_Wdata_ram : in std_logic_vector(31 downto 0) ;
  Min_data_ram_size : in std_logic_vector(5 downto 0) ;
  selector_IN_UNBOUNDED_acc_0_31017_31056 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31057 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31059 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31060 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31061 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31063 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31065 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31066 : in std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31068 : in std_logic;
  fuselector_MEMORY_CTRL_D21_251_i0_LOAD : in std_logic;
  fuselector_MEMORY_CTRL_D21_251_i0_STORE : in std_logic;
  selector_MUX_550_reg_13_0_0_0 : in std_logic;
  selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : in std_logic;
  selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : in std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : in std_logic;
  wrenable_reg_0 : in std_logic;
  wrenable_reg_1 : in std_logic;
  wrenable_reg_10 : in std_logic;
  wrenable_reg_11 : in std_logic;
  wrenable_reg_12 : in std_logic;
  wrenable_reg_13 : in std_logic;
  wrenable_reg_14 : in std_logic;
  wrenable_reg_15 : in std_logic;
  wrenable_reg_16 : in std_logic;
  wrenable_reg_17 : in std_logic;
  wrenable_reg_18 : in std_logic;
  wrenable_reg_19 : in std_logic;
  wrenable_reg_2 : in std_logic;
  wrenable_reg_20 : in std_logic;
  wrenable_reg_21 : in std_logic;
  wrenable_reg_22 : in std_logic;
  wrenable_reg_23 : in std_logic;
  wrenable_reg_24 : in std_logic;
  wrenable_reg_25 : in std_logic;
  wrenable_reg_26 : in std_logic;
  wrenable_reg_27 : in std_logic;
  wrenable_reg_28 : in std_logic;
  wrenable_reg_29 : in std_logic;
  wrenable_reg_3 : in std_logic;
  wrenable_reg_30 : in std_logic;
  wrenable_reg_31 : in std_logic;
  wrenable_reg_32 : in std_logic;
  wrenable_reg_33 : in std_logic;
  wrenable_reg_34 : in std_logic;
  wrenable_reg_35 : in std_logic;
  wrenable_reg_36 : in std_logic;
  wrenable_reg_37 : in std_logic;
  wrenable_reg_38 : in std_logic;
  wrenable_reg_39 : in std_logic;
  wrenable_reg_4 : in std_logic;
  wrenable_reg_40 : in std_logic;
  wrenable_reg_41 : in std_logic;
  wrenable_reg_42 : in std_logic;
  wrenable_reg_43 : in std_logic;
  wrenable_reg_44 : in std_logic;
  wrenable_reg_45 : in std_logic;
  wrenable_reg_46 : in std_logic;
  wrenable_reg_47 : in std_logic;
  wrenable_reg_5 : in std_logic;
  wrenable_reg_6 : in std_logic;
  wrenable_reg_7 : in std_logic;
  wrenable_reg_8 : in std_logic;
  wrenable_reg_9 : in std_logic;
  -- OUT
  Mout_oe_ram : out std_logic;
  Mout_we_ram : out std_logic;
  Mout_addr_ram : out std_logic_vector(31 downto 0) ;
  Mout_Wdata_ram : out std_logic_vector(31 downto 0) ;
  Mout_data_ram_size : out std_logic_vector(5 downto 0) ;
  OUT_MULTIIF_acc_0_31017_37300 : out std_logic_vector(0 downto 0);
  OUT_UNBOUNDED_acc_0_31017_31056 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31057 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31059 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31060 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31061 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31063 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31065 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31066 : out std_logic;
  OUT_UNBOUNDED_acc_0_31017_31068 : out std_logic

);
end datapath_acc_0;

architecture datapath_acc_0_arch of datapath_acc_0 is
  -- Component and signal declarations
  
  component constant_value
  generic(
   BITSIZE_out1: integer;
   value: std_logic_vector);
  port (
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component register_SE
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    wenable : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component register_STD
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    wenable : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component UUdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component extract_bit_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  
  component IUdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component lut_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in std_logic;
    in3 : in std_logic;
    in4 : in std_logic;
    in5 : in std_logic;
    in6 : in std_logic;
    in7 : in std_logic;
    in8 : in std_logic;
    in9 : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component UIdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component IIdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component multi_read_cond_FU
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component ui_extract_bit_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  
  component MEMORY_CTRL_D21
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_in3: integer;
   BITSIZE_out1: integer;
   BITSIZE_Min_addr_ram: integer;
   BITSIZE_Mout_addr_ram: integer;
   BITSIZE_M_Rdata_ram: integer;
   BITSIZE_Min_Wdata_ram: integer;
   BITSIZE_Mout_Wdata_ram: integer;
   BITSIZE_Min_data_ram_size: integer;
   BITSIZE_Mout_data_ram_size: integer);
  port (
    -- IN
    clock : in std_logic;
    start_port : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    in3 : in std_logic_vector(BITSIZE_in3-1 downto 0) ;
    in4 : in std_logic;
    sel_LOAD : in std_logic;
    sel_STORE : in std_logic;
    Min_oe_ram : in std_logic;
    Min_we_ram : in std_logic;
    Min_addr_ram : in std_logic_vector(BITSIZE_Min_addr_ram-1 downto 0) ;
    M_Rdata_ram : in std_logic_vector(BITSIZE_M_Rdata_ram-1 downto 0) ;
    Min_Wdata_ram : in std_logic_vector(BITSIZE_Min_Wdata_ram-1 downto 0) ;
    Min_data_ram_size : in std_logic_vector(BITSIZE_Min_data_ram_size-1 downto 0) ;
    M_DataRdy : in std_logic;
    -- OUT
    done_port : out std_logic;
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) ;
    Mout_oe_ram : out std_logic;
    Mout_we_ram : out std_logic;
    Mout_addr_ram : out std_logic_vector(BITSIZE_Mout_addr_ram-1 downto 0) ;
    Mout_Wdata_ram : out std_logic_vector(BITSIZE_Mout_Wdata_ram-1 downto 0) ;
    Mout_data_ram_size : out std_logic_vector(BITSIZE_Mout_data_ram_size-1 downto 0) 
  
  );
  end component;
  
  component bit_and_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component bit_ior_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component bit_not_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component eq_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component minus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component mult_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PIPE_PARAMETER: integer);
  port (
    -- IN
    clock : in std_logic;
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component negate_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component plus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_bit_and_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_bit_ior_concat_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_in3: integer;
   BITSIZE_out1: integer;
   OFFSET_PARAMETER: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    in3 : in unsigned (BITSIZE_in3-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_bit_ior_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_cond_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_in3: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    in3 : in unsigned (BITSIZE_in3-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_eq_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component ui_lshift_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PRECISION: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_mult_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PIPE_PARAMETER: integer);
  port (
    -- IN
    clock : in std_logic;
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_ne_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component ui_plus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_pointer_plus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   LSB_PARAMETER: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_rshift_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PRECISION: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_ternary_plus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_in3: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    in3 : in unsigned (BITSIZE_in3-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component bus_merger
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component OR_GATE
  generic(
   BITSIZE_in: integer;
   PORTSIZE_in: integer);
  port (
    -- IN
    \in\ : in std_logic_vector((PORTSIZE_in*BITSIZE_in)-1 downto 0) ;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  
  component ASSIGN_VECTOR_BOOL_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component MUX_GATE
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    sel : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  signal out_IIdata_converter_FU_111_i0_fu_acc_0_31017_37285 : signed (6 downto 0);
  signal out_IUdata_converter_FU_112_i0_fu_acc_0_31017_37291 : unsigned (7 downto 0);
  signal out_IUdata_converter_FU_15_i0_fu_acc_0_31017_36811 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_16_i0_fu_acc_0_31017_36817 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_250_i0_fu_acc_0_31017_37349 : unsigned (24 downto 0);
  signal out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_550_reg_13_0_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : std_logic_vector(31 downto 0) ;
  signal out_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : std_logic_vector(31 downto 0) ;
  signal out_UIdata_converter_FU_110_i0_fu_acc_0_31017_37279 : signed (5 downto 0);
  signal out_UIdata_converter_FU_161_i0_fu_acc_0_31017_37596 : signed (2 downto 0);
  signal out_UIdata_converter_FU_162_i0_fu_acc_0_31017_37599 : signed (1 downto 0);
  signal out_UIdata_converter_FU_165_i0_fu_acc_0_31017_37608 : signed (1 downto 0);
  signal out_UIdata_converter_FU_178_i0_fu_acc_0_31017_37668 : signed (2 downto 0);
  signal out_UIdata_converter_FU_179_i0_fu_acc_0_31017_37677 : signed (1 downto 0);
  signal out_UIdata_converter_FU_182_i0_fu_acc_0_31017_37689 : signed (1 downto 0);
  signal out_UIdata_converter_FU_189_i0_fu_acc_0_31017_37719 : signed (1 downto 0);
  signal out_UIdata_converter_FU_249_i0_fu_acc_0_31017_37343 : signed (1 downto 0);
  signal out_UUdata_converter_FU_109_i0_fu_acc_0_31017_37273 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_10_i0_fu_acc_0_31017_31597 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_113_i0_fu_acc_0_31017_31621 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_114_i0_fu_acc_0_31017_31629 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_117_i0_fu_acc_0_31017_33178 : std_logic_vector(30 downto 0) ;
  signal out_UUdata_converter_FU_118_i0_fu_acc_0_31017_33181 : std_logic_vector(30 downto 0) ;
  signal out_UUdata_converter_FU_119_i0_fu_acc_0_31017_37404 : std_logic_vector(7 downto 0) ;
  signal out_UUdata_converter_FU_11_i0_fu_acc_0_31017_31505 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_120_i0_fu_acc_0_31017_37417 : std_logic_vector(7 downto 0) ;
  signal out_UUdata_converter_FU_124_i0_fu_acc_0_31017_37434 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_12_i0_fu_acc_0_31017_31609 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_13_i0_fu_acc_0_31017_31518 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_149_i0_fu_acc_0_31017_37548 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_160_i0_fu_acc_0_31017_37584 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_164_i0_fu_acc_0_31017_37605 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_166_i0_fu_acc_0_31017_37617 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_177_i0_fu_acc_0_31017_37653 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_17_i0_fu_acc_0_31017_36820 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_181_i0_fu_acc_0_31017_37686 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_184_i0_fu_acc_0_31017_37701 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_185_i0_fu_acc_0_31017_37704 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_188_i0_fu_acc_0_31017_37716 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_190_i0_fu_acc_0_31017_37731 : std_logic_vector(9 downto 0) ;
  signal out_UUdata_converter_FU_195_i0_fu_acc_0_31017_37776 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_22_i0_fu_acc_0_31017_36907 : std_logic_vector(7 downto 0) ;
  signal out_UUdata_converter_FU_238_i0_fu_acc_0_31017_33175 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_23_i0_fu_acc_0_31017_36910 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_2_i0_fu_acc_0_31017_31544 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_3_i0_fu_acc_0_31017_31446 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_49_i0_fu_acc_0_31017_37015 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_4_i0_fu_acc_0_31017_31560 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_5_i0_fu_acc_0_31017_31466 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_62_i0_fu_acc_0_31017_37087 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_6_i0_fu_acc_0_31017_31573 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_7_i0_fu_acc_0_31017_31479 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_8_i0_fu_acc_0_31017_31585 : std_logic_vector(31 downto 0) ;
  signal out_UUdata_converter_FU_95_i0_fu_acc_0_31017_37222 : std_logic_vector(0 downto 0);
  signal out_UUdata_converter_FU_9_i0_fu_acc_0_31017_31492 : std_logic_vector(31 downto 0) ;
  signal out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674 : signed (1 downto 0);
  signal out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680 : signed (1 downto 0);
  signal out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692 : signed (1 downto 0);
  signal out_bit_ior_expr_FU_8_8_8_253_i0_fu_acc_0_31017_37671 : signed (2 downto 0);
  signal out_bit_not_expr_FU_8_8_254_i0_fu_acc_0_31017_37346 : signed (1 downto 0);
  signal out_const_0 : std_logic_vector(0 downto 0);
  signal out_const_1 : std_logic_vector(1 downto 0) ;
  signal out_const_10 : std_logic_vector(4 downto 0) ;
  signal out_const_11 : std_logic_vector(5 downto 0) ;
  signal out_const_12 : std_logic_vector(5 downto 0) ;
  signal out_const_13 : std_logic_vector(3 downto 0) ;
  signal out_const_14 : std_logic_vector(5 downto 0) ;
  signal out_const_15 : std_logic_vector(0 downto 0);
  signal out_const_16 : std_logic_vector(1 downto 0) ;
  signal out_const_17 : std_logic_vector(2 downto 0) ;
  signal out_const_18 : std_logic_vector(3 downto 0) ;
  signal out_const_19 : std_logic_vector(4 downto 0) ;
  signal out_const_2 : std_logic_vector(2 downto 0) ;
  signal out_const_20 : std_logic_vector(5 downto 0) ;
  signal out_const_21 : std_logic_vector(7 downto 0) ;
  signal out_const_22 : std_logic_vector(16 downto 0) ;
  signal out_const_23 : std_logic_vector(23 downto 0) ;
  signal out_const_24 : std_logic_vector(31 downto 0) ;
  signal out_const_25 : std_logic_vector(32 downto 0) ;
  signal out_const_26 : std_logic_vector(63 downto 0) ;
  signal out_const_27 : std_logic_vector(48 downto 0) ;
  signal out_const_28 : std_logic_vector(58 downto 0) ;
  signal out_const_29 : std_logic_vector(4 downto 0) ;
  signal out_const_3 : std_logic_vector(3 downto 0) ;
  signal out_const_30 : std_logic_vector(60 downto 0) ;
  signal out_const_31 : std_logic_vector(3 downto 0) ;
  signal out_const_32 : std_logic_vector(4 downto 0) ;
  signal out_const_33 : std_logic_vector(2 downto 0) ;
  signal out_const_34 : std_logic_vector(26 downto 0) ;
  signal out_const_35 : std_logic_vector(4 downto 0) ;
  signal out_const_36 : std_logic_vector(63 downto 0) ;
  signal out_const_37 : std_logic_vector(47 downto 0) ;
  signal out_const_38 : std_logic_vector(3 downto 0) ;
  signal out_const_39 : std_logic_vector(4 downto 0) ;
  signal out_const_4 : std_logic_vector(4 downto 0) ;
  signal out_const_40 : std_logic_vector(4 downto 0) ;
  signal out_const_41 : std_logic_vector(5 downto 0) ;
  signal out_const_42 : std_logic_vector(1 downto 0) ;
  signal out_const_43 : std_logic_vector(2 downto 0) ;
  signal out_const_44 : std_logic_vector(4 downto 0) ;
  signal out_const_45 : std_logic_vector(4 downto 0) ;
  signal out_const_46 : std_logic_vector(7 downto 0) ;
  signal out_const_47 : std_logic_vector(3 downto 0) ;
  signal out_const_48 : std_logic_vector(4 downto 0) ;
  signal out_const_49 : std_logic_vector(4 downto 0) ;
  signal out_const_5 : std_logic_vector(5 downto 0) ;
  signal out_const_50 : std_logic_vector(7 downto 0) ;
  signal out_const_51 : std_logic_vector(2 downto 0) ;
  signal out_const_52 : std_logic_vector(4 downto 0) ;
  signal out_const_53 : std_logic_vector(7 downto 0) ;
  signal out_const_54 : std_logic_vector(55 downto 0) ;
  signal out_const_55 : std_logic_vector(11 downto 0) ;
  signal out_const_56 : std_logic_vector(10 downto 0) ;
  signal out_const_57 : std_logic_vector(4 downto 0) ;
  signal out_const_58 : std_logic_vector(7 downto 0) ;
  signal out_const_59 : std_logic_vector(3 downto 0) ;
  signal out_const_6 : std_logic_vector(6 downto 0) ;
  signal out_const_60 : std_logic_vector(4 downto 0) ;
  signal out_const_61 : std_logic_vector(31 downto 0) ;
  signal out_const_62 : std_logic_vector(4 downto 0) ;
  signal out_const_63 : std_logic_vector(31 downto 0) ;
  signal out_const_64 : std_logic_vector(5 downto 0) ;
  signal out_const_65 : std_logic_vector(7 downto 0) ;
  signal out_const_66 : std_logic_vector(30 downto 0) ;
  signal out_const_67 : std_logic_vector(9 downto 0) ;
  signal out_const_68 : std_logic_vector(47 downto 0) ;
  signal out_const_69 : std_logic_vector(63 downto 0) ;
  signal out_const_7 : std_logic_vector(8 downto 0) ;
  signal out_const_70 : std_logic_vector(16 downto 0) ;
  signal out_const_71 : std_logic_vector(16 downto 0) ;
  signal out_const_72 : std_logic_vector(31 downto 0) ;
  signal out_const_73 : std_logic_vector(22 downto 0) ;
  signal out_const_74 : std_logic_vector(31 downto 0) ;
  signal out_const_75 : std_logic_vector(30 downto 0) ;
  signal out_const_76 : std_logic_vector(31 downto 0) ;
  signal out_const_77 : std_logic_vector(32 downto 0) ;
  signal out_const_78 : std_logic_vector(46 downto 0) ;
  signal out_const_8 : std_logic_vector(5 downto 0) ;
  signal out_const_9 : std_logic_vector(5 downto 0) ;
  signal out_conv_out_const_6_7_6 : std_logic_vector(5 downto 0) ;
  signal out_eq_expr_FU_32_0_32_255_i0_fu_acc_0_31017_36800 : std_logic_vector(0 downto 0);
  signal out_eq_expr_FU_32_0_32_256_i0_fu_acc_0_31017_36808 : std_logic_vector(0 downto 0);
  signal out_extract_bit_expr_FU_14_i0_fu_acc_0_31017_36805 : std_logic;
  signal out_extract_bit_expr_FU_18_i0_fu_acc_0_31017_36832 : std_logic;
  signal out_extract_bit_expr_FU_198_i0_fu_acc_0_31017_37788 : std_logic;
  signal out_extract_bit_expr_FU_199_i0_fu_acc_0_31017_37791 : std_logic;
  signal out_extract_bit_expr_FU_201_i0_fu_acc_0_31017_37797 : std_logic;
  signal out_extract_bit_expr_FU_213_i0_fu_acc_0_31017_37839 : std_logic;
  signal out_extract_bit_expr_FU_214_i0_fu_acc_0_31017_37842 : std_logic;
  signal out_extract_bit_expr_FU_216_i0_fu_acc_0_31017_37848 : std_logic;
  signal out_extract_bit_expr_FU_218_i0_fu_acc_0_31017_37854 : std_logic;
  signal out_extract_bit_expr_FU_219_i0_fu_acc_0_31017_37857 : std_logic;
  signal out_extract_bit_expr_FU_221_i0_fu_acc_0_31017_37863 : std_logic;
  signal out_extract_bit_expr_FU_227_i0_fu_acc_0_31017_37881 : std_logic;
  signal out_extract_bit_expr_FU_228_i0_fu_acc_0_31017_37884 : std_logic;
  signal out_extract_bit_expr_FU_230_i0_fu_acc_0_31017_37890 : std_logic;
  signal out_extract_bit_expr_FU_233_i0_fu_acc_0_31017_37914 : std_logic;
  signal out_extract_bit_expr_FU_234_i0_fu_acc_0_31017_37917 : std_logic;
  signal out_extract_bit_expr_FU_236_i0_fu_acc_0_31017_37923 : std_logic;
  signal out_extract_bit_expr_FU_26_i0_fu_acc_0_31017_36943 : std_logic;
  signal out_extract_bit_expr_FU_27_i0_fu_acc_0_31017_36946 : std_logic;
  signal out_extract_bit_expr_FU_28_i0_fu_acc_0_31017_36949 : std_logic;
  signal out_extract_bit_expr_FU_29_i0_fu_acc_0_31017_36952 : std_logic;
  signal out_extract_bit_expr_FU_30_i0_fu_acc_0_31017_36955 : std_logic;
  signal out_extract_bit_expr_FU_31_i0_fu_acc_0_31017_36958 : std_logic;
  signal out_extract_bit_expr_FU_32_i0_fu_acc_0_31017_36961 : std_logic;
  signal out_extract_bit_expr_FU_33_i0_fu_acc_0_31017_36964 : std_logic;
  signal out_extract_bit_expr_FU_34_i0_fu_acc_0_31017_36967 : std_logic;
  signal out_extract_bit_expr_FU_35_i0_fu_acc_0_31017_36970 : std_logic;
  signal out_extract_bit_expr_FU_36_i0_fu_acc_0_31017_36973 : std_logic;
  signal out_extract_bit_expr_FU_37_i0_fu_acc_0_31017_36976 : std_logic;
  signal out_extract_bit_expr_FU_38_i0_fu_acc_0_31017_36979 : std_logic;
  signal out_extract_bit_expr_FU_39_i0_fu_acc_0_31017_36982 : std_logic;
  signal out_extract_bit_expr_FU_40_i0_fu_acc_0_31017_36985 : std_logic;
  signal out_extract_bit_expr_FU_41_i0_fu_acc_0_31017_36988 : std_logic;
  signal out_extract_bit_expr_FU_50_i0_fu_acc_0_31017_37021 : std_logic;
  signal out_extract_bit_expr_FU_51_i0_fu_acc_0_31017_37024 : std_logic;
  signal out_extract_bit_expr_FU_52_i0_fu_acc_0_31017_37027 : std_logic;
  signal out_extract_bit_expr_FU_53_i0_fu_acc_0_31017_37030 : std_logic;
  signal out_extract_bit_expr_FU_54_i0_fu_acc_0_31017_37033 : std_logic;
  signal out_extract_bit_expr_FU_55_i0_fu_acc_0_31017_37036 : std_logic;
  signal out_extract_bit_expr_FU_56_i0_fu_acc_0_31017_37039 : std_logic;
  signal out_extract_bit_expr_FU_57_i0_fu_acc_0_31017_37042 : std_logic;
  signal out_extract_bit_expr_FU_63_i0_fu_acc_0_31017_37126 : std_logic;
  signal out_extract_bit_expr_FU_64_i0_fu_acc_0_31017_37129 : std_logic;
  signal out_extract_bit_expr_FU_65_i0_fu_acc_0_31017_37132 : std_logic;
  signal out_extract_bit_expr_FU_66_i0_fu_acc_0_31017_37135 : std_logic;
  signal out_extract_bit_expr_FU_67_i0_fu_acc_0_31017_37138 : std_logic;
  signal out_extract_bit_expr_FU_68_i0_fu_acc_0_31017_37141 : std_logic;
  signal out_extract_bit_expr_FU_69_i0_fu_acc_0_31017_37144 : std_logic;
  signal out_extract_bit_expr_FU_70_i0_fu_acc_0_31017_37147 : std_logic;
  signal out_extract_bit_expr_FU_71_i0_fu_acc_0_31017_37150 : std_logic;
  signal out_extract_bit_expr_FU_72_i0_fu_acc_0_31017_37153 : std_logic;
  signal out_extract_bit_expr_FU_73_i0_fu_acc_0_31017_37156 : std_logic;
  signal out_extract_bit_expr_FU_74_i0_fu_acc_0_31017_37159 : std_logic;
  signal out_extract_bit_expr_FU_75_i0_fu_acc_0_31017_37162 : std_logic;
  signal out_extract_bit_expr_FU_76_i0_fu_acc_0_31017_37165 : std_logic;
  signal out_extract_bit_expr_FU_77_i0_fu_acc_0_31017_37168 : std_logic;
  signal out_extract_bit_expr_FU_78_i0_fu_acc_0_31017_37171 : std_logic;
  signal out_extract_bit_expr_FU_79_i0_fu_acc_0_31017_37174 : std_logic;
  signal out_extract_bit_expr_FU_80_i0_fu_acc_0_31017_37177 : std_logic;
  signal out_extract_bit_expr_FU_81_i0_fu_acc_0_31017_37180 : std_logic;
  signal out_extract_bit_expr_FU_82_i0_fu_acc_0_31017_37183 : std_logic;
  signal out_extract_bit_expr_FU_83_i0_fu_acc_0_31017_37186 : std_logic;
  signal out_extract_bit_expr_FU_84_i0_fu_acc_0_31017_37189 : std_logic;
  signal out_extract_bit_expr_FU_85_i0_fu_acc_0_31017_37192 : std_logic;
  signal out_extract_bit_expr_FU_86_i0_fu_acc_0_31017_37195 : std_logic;
  signal out_extract_bit_expr_FU_87_i0_fu_acc_0_31017_37198 : std_logic;
  signal out_extract_bit_expr_FU_88_i0_fu_acc_0_31017_37201 : std_logic;
  signal out_extract_bit_expr_FU_89_i0_fu_acc_0_31017_37204 : std_logic;
  signal out_extract_bit_expr_FU_90_i0_fu_acc_0_31017_37207 : std_logic;
  signal out_extract_bit_expr_FU_91_i0_fu_acc_0_31017_37210 : std_logic;
  signal out_extract_bit_expr_FU_92_i0_fu_acc_0_31017_37213 : std_logic;
  signal out_extract_bit_expr_FU_93_i0_fu_acc_0_31017_37216 : std_logic;
  signal out_extract_bit_expr_FU_94_i0_fu_acc_0_31017_37219 : std_logic;
  signal out_iu_conv_conn_obj_0_IUdata_converter_FU_iu_conv_0 : unsigned (31 downto 0);
  signal out_iu_conv_conn_obj_1_IUdata_converter_FU_iu_conv_1 : unsigned (31 downto 0);
  signal out_lut_expr_FU_100_i0_fu_acc_0_31017_37246 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_101_i0_fu_acc_0_31017_37249 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_102_i0_fu_acc_0_31017_37252 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_103_i0_fu_acc_0_31017_37255 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_104_i0_fu_acc_0_31017_37258 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_105_i0_fu_acc_0_31017_37261 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_106_i0_fu_acc_0_31017_37264 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_107_i0_fu_acc_0_31017_37267 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_108_i0_fu_acc_0_31017_37270 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_123_i0_fu_acc_0_31017_37431 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_133_i0_fu_acc_0_31017_38089 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_134_i0_fu_acc_0_31017_38092 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_135_i0_fu_acc_0_31017_37473 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_136_i0_fu_acc_0_31017_37479 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_145_i0_fu_acc_0_31017_38097 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_146_i0_fu_acc_0_31017_38100 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_147_i0_fu_acc_0_31017_37518 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_148_i0_fu_acc_0_31017_37524 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_158_i0_fu_acc_0_31017_38105 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_159_i0_fu_acc_0_31017_37581 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_163_i0_fu_acc_0_31017_37602 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_175_i0_fu_acc_0_31017_38110 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_176_i0_fu_acc_0_31017_37650 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_180_i0_fu_acc_0_31017_37683 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_187_i0_fu_acc_0_31017_37713 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_194_i0_fu_acc_0_31017_37773 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_19_i0_fu_acc_0_31017_36835 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_202_i0_fu_acc_0_31017_38117 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_203_i0_fu_acc_0_31017_37803 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_20_i0_fu_acc_0_31017_36838 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_217_i0_fu_acc_0_31017_37851 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_222_i0_fu_acc_0_31017_38122 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_223_i0_fu_acc_0_31017_38125 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_224_i0_fu_acc_0_31017_38128 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_225_i0_fu_acc_0_31017_38132 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_226_i0_fu_acc_0_31017_37878 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_231_i0_fu_acc_0_31017_38137 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_232_i0_fu_acc_0_31017_37896 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_237_i0_fu_acc_0_31017_37926 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_247_i0_fu_acc_0_31017_37337 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_248_i0_fu_acc_0_31017_37340 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_24_i0_fu_acc_0_31017_36916 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_25_i0_fu_acc_0_31017_36919 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_42_i0_fu_acc_0_31017_36991 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_43_i0_fu_acc_0_31017_36994 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_44_i0_fu_acc_0_31017_36997 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_45_i0_fu_acc_0_31017_37000 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_46_i0_fu_acc_0_31017_37003 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_47_i0_fu_acc_0_31017_37009 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_48_i0_fu_acc_0_31017_37012 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_58_i0_fu_acc_0_31017_37045 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_59_i0_fu_acc_0_31017_37048 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_60_i0_fu_acc_0_31017_37051 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_61_i0_fu_acc_0_31017_37054 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_96_i0_fu_acc_0_31017_37234 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_97_i0_fu_acc_0_31017_37237 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_98_i0_fu_acc_0_31017_37240 : std_logic_vector(0 downto 0);
  signal out_lut_expr_FU_99_i0_fu_acc_0_31017_37243 : std_logic_vector(0 downto 0);
  signal out_minus_expr_FU_0_8_8_257_i0_fu_acc_0_31017_37288 : signed (8 downto 0);
  signal out_mult_expr_FU_32_32_32_0_258_i0_fu_acc_0_31017_31062 : signed (31 downto 0);
  signal out_multi_read_cond_FU_115_i0_fu_acc_0_31017_37300 : std_logic_vector(0 downto 0);
  signal out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814 : signed (31 downto 0);
  signal out_plus_expr_FU_32_32_32_260_i0_fu_acc_0_31017_31058 : signed (31 downto 0);
  signal out_plus_expr_FU_8_0_8_261_i0_fu_acc_0_31017_37282 : signed (6 downto 0);
  signal out_reg_0_reg_0 : std_logic_vector(31 downto 0) ;
  signal out_reg_10_reg_10 : std_logic_vector(31 downto 0) ;
  signal out_reg_11_reg_11 : std_logic_vector(31 downto 0) ;
  signal out_reg_12_reg_12 : std_logic_vector(0 downto 0);
  signal out_reg_13_reg_13 : std_logic_vector(31 downto 0) ;
  signal out_reg_14_reg_14 : std_logic_vector(31 downto 0) ;
  signal out_reg_15_reg_15 : std_logic_vector(6 downto 0) ;
  signal out_reg_16_reg_16 : std_logic_vector(7 downto 0) ;
  signal out_reg_17_reg_17 : std_logic_vector(31 downto 0) ;
  signal out_reg_18_reg_18 : std_logic_vector(31 downto 0) ;
  signal out_reg_19_reg_19 : std_logic_vector(31 downto 0) ;
  signal out_reg_1_reg_1 : std_logic_vector(31 downto 0) ;
  signal out_reg_20_reg_20 : std_logic_vector(7 downto 0) ;
  signal out_reg_21_reg_21 : std_logic_vector(0 downto 0);
  signal out_reg_22_reg_22 : std_logic_vector(0 downto 0);
  signal out_reg_23_reg_23 : std_logic_vector(23 downto 0) ;
  signal out_reg_24_reg_24 : std_logic_vector(2 downto 0) ;
  signal out_reg_25_reg_25 : std_logic_vector(1 downto 0) ;
  signal out_reg_26_reg_26 : std_logic_vector(1 downto 0) ;
  signal out_reg_27_reg_27 : std_logic_vector(0 downto 0);
  signal out_reg_28_reg_28 : std_logic_vector(0 downto 0);
  signal out_reg_29_reg_29 : std_logic_vector(31 downto 0) ;
  signal out_reg_2_reg_2 : std_logic_vector(31 downto 0) ;
  signal out_reg_30_reg_30 : std_logic_vector(31 downto 0) ;
  signal out_reg_31_reg_31 : std_logic_vector(31 downto 0) ;
  signal out_reg_32_reg_32 : std_logic_vector(9 downto 0) ;
  signal out_reg_33_reg_33 : std_logic_vector(47 downto 0) ;
  signal out_reg_34_reg_34 : std_logic_vector(0 downto 0);
  signal out_reg_35_reg_35 : std_logic_vector(1 downto 0) ;
  signal out_reg_36_reg_36 : std_logic_vector(0 downto 0);
  signal out_reg_37_reg_37 : std_logic_vector(0 downto 0);
  signal out_reg_38_reg_38 : std_logic_vector(0 downto 0);
  signal out_reg_39_reg_39 : std_logic_vector(0 downto 0);
  signal out_reg_3_reg_3 : std_logic_vector(31 downto 0) ;
  signal out_reg_40_reg_40 : std_logic_vector(0 downto 0);
  signal out_reg_41_reg_41 : std_logic_vector(0 downto 0);
  signal out_reg_42_reg_42 : std_logic_vector(0 downto 0);
  signal out_reg_43_reg_43 : std_logic_vector(0 downto 0);
  signal out_reg_44_reg_44 : std_logic_vector(0 downto 0);
  signal out_reg_45_reg_45 : std_logic_vector(31 downto 0) ;
  signal out_reg_46_reg_46 : std_logic_vector(0 downto 0);
  signal out_reg_47_reg_47 : std_logic_vector(31 downto 0) ;
  signal out_reg_4_reg_4 : std_logic_vector(31 downto 0) ;
  signal out_reg_5_reg_5 : std_logic_vector(31 downto 0) ;
  signal out_reg_6_reg_6 : std_logic_vector(31 downto 0) ;
  signal out_reg_7_reg_7 : std_logic_vector(31 downto 0) ;
  signal out_reg_8_reg_8 : std_logic_vector(31 downto 0) ;
  signal out_reg_9_reg_9 : std_logic_vector(31 downto 0) ;
  signal out_ui_bit_and_expr_FU_0_32_32_262_i0_fu_acc_0_31017_37833 : unsigned (30 downto 0);
  signal out_ui_bit_and_expr_FU_0_64_64_263_i0_fu_acc_0_31017_37725 : unsigned (46 downto 0);
  signal out_ui_bit_and_expr_FU_0_64_64_264_i0_fu_acc_0_31017_37746 : unsigned (32 downto 0);
  signal out_ui_bit_and_expr_FU_0_8_8_265_i0_fu_acc_0_31017_37414 : unsigned (7 downto 0);
  signal out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665 : unsigned (0 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_267_i0_fu_acc_0_31017_37358 : unsigned (24 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_268_i0_fu_acc_0_31017_37367 : unsigned (22 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_269_i0_fu_acc_0_31017_37393 : unsigned (22 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_269_i1_fu_acc_0_31017_37422 : unsigned (22 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_269_i2_fu_acc_0_31017_37740 : unsigned (22 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_269_i3_fu_acc_0_31017_37755 : unsigned (22 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_270_i0_fu_acc_0_31017_37536 : unsigned (23 downto 0);
  signal out_ui_bit_and_expr_FU_32_0_32_270_i1_fu_acc_0_31017_37539 : unsigned (23 downto 0);
  signal out_ui_bit_and_expr_FU_32_32_32_271_i0_fu_acc_0_31017_37352 : unsigned (24 downto 0);
  signal out_ui_bit_and_expr_FU_8_0_8_272_i0_fu_acc_0_31017_36877 : unsigned (5 downto 0);
  signal out_ui_bit_and_expr_FU_8_0_8_273_i0_fu_acc_0_31017_36904 : unsigned (7 downto 0);
  signal out_ui_bit_and_expr_FU_8_0_8_274_i0_fu_acc_0_31017_37078 : unsigned (1 downto 0);
  signal out_ui_bit_and_expr_FU_8_0_8_275_i0_fu_acc_0_31017_37401 : unsigned (7 downto 0);
  signal out_ui_bit_ior_concat_expr_FU_276_i0_fu_acc_0_31017_37361 : unsigned (31 downto 0);
  signal out_ui_bit_ior_concat_expr_FU_277_i0_fu_acc_0_31017_37385 : unsigned (31 downto 0);
  signal out_ui_bit_ior_expr_FU_0_32_32_278_i0_fu_acc_0_31017_37530 : unsigned (23 downto 0);
  signal out_ui_bit_ior_expr_FU_0_32_32_278_i1_fu_acc_0_31017_37533 : unsigned (23 downto 0);
  signal out_ui_bit_ior_expr_FU_0_32_32_279_i0_fu_acc_0_31017_37542 : unsigned (31 downto 0);
  signal out_ui_bit_ior_expr_FU_0_32_32_280_i0_fu_acc_0_31017_37836 : unsigned (31 downto 0);
  signal out_ui_bit_ior_expr_FU_0_64_64_281_i0_fu_acc_0_31017_37743 : unsigned (32 downto 0);
  signal out_ui_bit_ior_expr_FU_0_8_8_282_i0_fu_acc_0_31017_37093 : unsigned (4 downto 0);
  signal out_ui_bit_ior_expr_FU_0_8_8_283_i0_fu_acc_0_31017_37228 : unsigned (2 downto 0);
  signal out_ui_bit_ior_expr_FU_0_8_8_284_i0_fu_acc_0_31017_37231 : unsigned (4 downto 0);
  signal out_ui_bit_ior_expr_FU_0_8_8_285_i0_fu_acc_0_31017_37276 : unsigned (4 downto 0);
  signal out_ui_bit_ior_expr_FU_8_8_8_286_i0_fu_acc_0_31017_37587 : unsigned (1 downto 0);
  signal out_ui_bit_ior_expr_FU_8_8_8_286_i1_fu_acc_0_31017_37590 : unsigned (1 downto 0);
  signal out_ui_bit_ior_expr_FU_8_8_8_286_i2_fu_acc_0_31017_37656 : unsigned (1 downto 0);
  signal out_ui_bit_ior_expr_FU_8_8_8_286_i3_fu_acc_0_31017_37659 : unsigned (1 downto 0);
  signal out_ui_cond_expr_FU_16_16_16_16_287_i0_fu_acc_0_31017_37908 : unsigned (9 downto 0);
  signal out_ui_cond_expr_FU_16_16_16_16_287_i1_fu_acc_0_31017_37935 : unsigned (9 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i0_fu_acc_0_31017_36847 : unsigned (31 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i1_fu_acc_0_31017_37006 : unsigned (23 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i2_fu_acc_0_31017_37063 : unsigned (21 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i3_fu_acc_0_31017_37108 : unsigned (17 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i4_fu_acc_0_31017_37899 : unsigned (31 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i5_fu_acc_0_31017_37902 : unsigned (31 downto 0);
  signal out_ui_cond_expr_FU_32_32_32_32_288_i6_fu_acc_0_31017_37941 : unsigned (31 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i0_fu_acc_0_31017_36841 : unsigned (7 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i1_fu_acc_0_31017_36934 : unsigned (5 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i2_fu_acc_0_31017_37370 : unsigned (7 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i3_fu_acc_0_31017_37482 : unsigned (1 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i4_fu_acc_0_31017_37527 : unsigned (1 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i5_fu_acc_0_31017_37545 : unsigned (1 downto 0);
  signal out_ui_cond_expr_FU_8_8_8_8_289_i6_fu_acc_0_31017_37614 : unsigned (1 downto 0);
  signal out_ui_eq_expr_FU_16_0_16_290_i0_fu_acc_0_31017_36856 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_16_0_16_290_i2_fu_acc_0_31017_36868 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i1_fu_acc_0_31017_36895 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i2_fu_acc_0_31017_36901 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i3_fu_acc_0_31017_37120 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i4_fu_acc_0_31017_37123 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_292_i0_fu_acc_0_31017_37355 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_293_i0_fu_acc_0_31017_37440 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_293_i1_fu_acc_0_31017_37485 : std_logic_vector(0 downto 0);
  signal out_ui_extract_bit_expr_FU_121_i0_fu_acc_0_31017_37951 : std_logic;
  signal out_ui_extract_bit_expr_FU_122_i0_fu_acc_0_31017_37955 : std_logic;
  signal out_ui_extract_bit_expr_FU_125_i0_fu_acc_0_31017_37959 : std_logic;
  signal out_ui_extract_bit_expr_FU_126_i0_fu_acc_0_31017_37963 : std_logic;
  signal out_ui_extract_bit_expr_FU_127_i0_fu_acc_0_31017_37967 : std_logic;
  signal out_ui_extract_bit_expr_FU_128_i0_fu_acc_0_31017_37971 : std_logic;
  signal out_ui_extract_bit_expr_FU_129_i0_fu_acc_0_31017_37975 : std_logic;
  signal out_ui_extract_bit_expr_FU_130_i0_fu_acc_0_31017_37979 : std_logic;
  signal out_ui_extract_bit_expr_FU_131_i0_fu_acc_0_31017_37983 : std_logic;
  signal out_ui_extract_bit_expr_FU_132_i0_fu_acc_0_31017_37987 : std_logic;
  signal out_ui_extract_bit_expr_FU_137_i0_fu_acc_0_31017_37991 : std_logic;
  signal out_ui_extract_bit_expr_FU_138_i0_fu_acc_0_31017_37995 : std_logic;
  signal out_ui_extract_bit_expr_FU_139_i0_fu_acc_0_31017_37999 : std_logic;
  signal out_ui_extract_bit_expr_FU_140_i0_fu_acc_0_31017_38003 : std_logic;
  signal out_ui_extract_bit_expr_FU_141_i0_fu_acc_0_31017_38007 : std_logic;
  signal out_ui_extract_bit_expr_FU_142_i0_fu_acc_0_31017_38011 : std_logic;
  signal out_ui_extract_bit_expr_FU_143_i0_fu_acc_0_31017_38015 : std_logic;
  signal out_ui_extract_bit_expr_FU_144_i0_fu_acc_0_31017_38019 : std_logic;
  signal out_ui_extract_bit_expr_FU_150_i0_fu_acc_0_31017_38023 : std_logic;
  signal out_ui_extract_bit_expr_FU_151_i0_fu_acc_0_31017_38027 : std_logic;
  signal out_ui_extract_bit_expr_FU_152_i0_fu_acc_0_31017_38031 : std_logic;
  signal out_ui_extract_bit_expr_FU_153_i0_fu_acc_0_31017_38035 : std_logic;
  signal out_ui_extract_bit_expr_FU_154_i0_fu_acc_0_31017_38039 : std_logic;
  signal out_ui_extract_bit_expr_FU_155_i0_fu_acc_0_31017_38043 : std_logic;
  signal out_ui_extract_bit_expr_FU_156_i0_fu_acc_0_31017_38047 : std_logic;
  signal out_ui_extract_bit_expr_FU_157_i0_fu_acc_0_31017_38051 : std_logic;
  signal out_ui_extract_bit_expr_FU_167_i0_fu_acc_0_31017_38055 : std_logic;
  signal out_ui_extract_bit_expr_FU_168_i0_fu_acc_0_31017_38059 : std_logic;
  signal out_ui_extract_bit_expr_FU_169_i0_fu_acc_0_31017_38063 : std_logic;
  signal out_ui_extract_bit_expr_FU_170_i0_fu_acc_0_31017_38067 : std_logic;
  signal out_ui_extract_bit_expr_FU_171_i0_fu_acc_0_31017_38071 : std_logic;
  signal out_ui_extract_bit_expr_FU_172_i0_fu_acc_0_31017_38075 : std_logic;
  signal out_ui_extract_bit_expr_FU_173_i0_fu_acc_0_31017_38079 : std_logic;
  signal out_ui_extract_bit_expr_FU_174_i0_fu_acc_0_31017_38083 : std_logic;
  signal out_ui_extract_bit_expr_FU_183_i0_fu_acc_0_31017_37698 : std_logic;
  signal out_ui_extract_bit_expr_FU_186_i0_fu_acc_0_31017_37710 : std_logic;
  signal out_ui_extract_bit_expr_FU_191_i0_fu_acc_0_31017_37749 : std_logic;
  signal out_ui_extract_bit_expr_FU_192_i0_fu_acc_0_31017_37767 : std_logic;
  signal out_ui_extract_bit_expr_FU_193_i0_fu_acc_0_31017_37770 : std_logic;
  signal out_ui_extract_bit_expr_FU_196_i0_fu_acc_0_31017_37782 : std_logic;
  signal out_ui_extract_bit_expr_FU_197_i0_fu_acc_0_31017_37785 : std_logic;
  signal out_ui_extract_bit_expr_FU_200_i0_fu_acc_0_31017_37794 : std_logic;
  signal out_ui_extract_bit_expr_FU_204_i0_fu_acc_0_31017_37806 : std_logic;
  signal out_ui_extract_bit_expr_FU_205_i0_fu_acc_0_31017_37809 : std_logic;
  signal out_ui_extract_bit_expr_FU_206_i0_fu_acc_0_31017_37812 : std_logic;
  signal out_ui_extract_bit_expr_FU_207_i0_fu_acc_0_31017_37815 : std_logic;
  signal out_ui_extract_bit_expr_FU_208_i0_fu_acc_0_31017_37818 : std_logic;
  signal out_ui_extract_bit_expr_FU_209_i0_fu_acc_0_31017_37821 : std_logic;
  signal out_ui_extract_bit_expr_FU_210_i0_fu_acc_0_31017_37824 : std_logic;
  signal out_ui_extract_bit_expr_FU_211_i0_fu_acc_0_31017_37827 : std_logic;
  signal out_ui_extract_bit_expr_FU_212_i0_fu_acc_0_31017_37830 : std_logic;
  signal out_ui_extract_bit_expr_FU_215_i0_fu_acc_0_31017_37845 : std_logic;
  signal out_ui_extract_bit_expr_FU_220_i0_fu_acc_0_31017_37860 : std_logic;
  signal out_ui_extract_bit_expr_FU_229_i0_fu_acc_0_31017_37887 : std_logic;
  signal out_ui_extract_bit_expr_FU_235_i0_fu_acc_0_31017_37920 : std_logic;
  signal out_ui_extract_bit_expr_FU_240_i0_fu_acc_0_31017_37316 : std_logic;
  signal out_ui_extract_bit_expr_FU_241_i0_fu_acc_0_31017_37319 : std_logic;
  signal out_ui_extract_bit_expr_FU_242_i0_fu_acc_0_31017_37322 : std_logic;
  signal out_ui_extract_bit_expr_FU_243_i0_fu_acc_0_31017_37325 : std_logic;
  signal out_ui_extract_bit_expr_FU_244_i0_fu_acc_0_31017_37328 : std_logic;
  signal out_ui_extract_bit_expr_FU_245_i0_fu_acc_0_31017_37331 : std_logic;
  signal out_ui_extract_bit_expr_FU_246_i0_fu_acc_0_31017_37334 : std_logic;
  signal out_ui_lshift_expr_FU_32_0_32_294_i0_fu_acc_0_31017_36823 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_294_i1_fu_acc_0_31017_37437 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_295_i0_fu_acc_0_31017_36829 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_296_i0_fu_acc_0_31017_36844 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_297_i0_fu_acc_0_31017_37066 : unsigned (23 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_298_i0_fu_acc_0_31017_37111 : unsigned (18 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_298_i1_fu_acc_0_31017_37114 : unsigned (19 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_298_i2_fu_acc_0_31017_37758 : unsigned (23 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_299_i0_fu_acc_0_31017_37294 : unsigned (30 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_300_i0_fu_acc_0_31017_37310 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_301_i0_fu_acc_0_31017_37373 : unsigned (30 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_301_i1_fu_acc_0_31017_37382 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_302_i0_fu_acc_0_31017_37911 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_0_32_302_i1_fu_acc_0_31017_37938 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301 : unsigned (31 downto 0);
  signal out_ui_lshift_expr_FU_64_0_64_304_i0_fu_acc_0_31017_37728 : unsigned (47 downto 0);
  signal out_ui_lshift_expr_FU_64_0_64_305_i0_fu_acc_0_31017_37734 : unsigned (32 downto 0);
  signal out_ui_lshift_expr_FU_64_64_64_306_i0_fu_acc_0_31017_37722 : unsigned (46 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i0_fu_acc_0_31017_36880 : unsigned (6 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i1_fu_acc_0_31017_36883 : unsigned (7 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i2_fu_acc_0_31017_36937 : unsigned (6 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i3_fu_acc_0_31017_36940 : unsigned (7 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i4_fu_acc_0_31017_37081 : unsigned (2 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_307_i5_fu_acc_0_31017_37084 : unsigned (3 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_308_i0_fu_acc_0_31017_36913 : unsigned (4 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_309_i0_fu_acc_0_31017_37018 : unsigned (3 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_310_i0_fu_acc_0_31017_37090 : unsigned (2 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_311_i0_fu_acc_0_31017_37225 : unsigned (1 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_312_i0_fu_acc_0_31017_37551 : unsigned (1 downto 0);
  signal out_ui_lshift_expr_FU_8_0_8_312_i1_fu_acc_0_31017_37620 : unsigned (1 downto 0);
  signal out_ui_mult_expr_FU_32_32_32_0_313_i0_fu_acc_0_31017_37695 : unsigned (47 downto 0);
  signal out_ui_ne_expr_FU_32_0_32_314_i0_fu_acc_0_31017_37476 : std_logic_vector(0 downto 0);
  signal out_ui_ne_expr_FU_32_0_32_314_i1_fu_acc_0_31017_37521 : std_logic_vector(0 downto 0);
  signal out_ui_ne_expr_FU_32_0_32_315_i0_fu_acc_0_31017_37764 : std_logic_vector(0 downto 0);
  signal out_ui_plus_expr_FU_0_32_32_316_i0_fu_acc_0_31017_37307 : unsigned (25 downto 0);
  signal out_ui_plus_expr_FU_16_16_16_317_i0_fu_acc_0_31017_37707 : unsigned (9 downto 0);
  signal out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779 : unsigned (32 downto 0);
  signal out_ui_plus_expr_FU_8_8_8_319_i0_fu_acc_0_31017_37379 : unsigned (8 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_320_i0_fu_acc_0_31017_31501 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_320_i1_fu_acc_0_31017_31514 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_320_i2_fu_acc_0_31017_31527 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_321_i0_fu_acc_0_31017_31564 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_321_i1_fu_acc_0_31017_31600 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_321_i2_fu_acc_0_31017_31632 : unsigned (31 downto 0);
  signal out_ui_pointer_plus_expr_FU_32_0_32_322_i0_fu_acc_0_31017_31625 : unsigned (31 downto 0);
  signal out_ui_rshift_expr_FU_16_0_16_323_i0_fu_acc_0_31017_36871 : unsigned (6 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_324_i0_fu_acc_0_31017_36826 : unsigned (0 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_325_i0_fu_acc_0_31017_36853 : unsigned (15 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_326_i0_fu_acc_0_31017_36862 : unsigned (7 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_327_i0_fu_acc_0_31017_36865 : unsigned (11 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_328_i0_fu_acc_0_31017_36886 : unsigned (23 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_329_i0_fu_acc_0_31017_36892 : unsigned (19 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_330_i0_fu_acc_0_31017_36898 : unsigned (27 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_330_i1_fu_acc_0_31017_37069 : unsigned (19 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_331_i0_fu_acc_0_31017_37057 : unsigned (21 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_332_i0_fu_acc_0_31017_37072 : unsigned (2 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_332_i1_fu_acc_0_31017_37099 : unsigned (18 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_332_i2_fu_acc_0_31017_37105 : unsigned (17 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_332_i3_fu_acc_0_31017_37761 : unsigned (22 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_333_i0_fu_acc_0_31017_37117 : unsigned (17 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_334_i0_fu_acc_0_31017_37297 : unsigned (7 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_334_i1_fu_acc_0_31017_37364 : unsigned (8 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_334_i2_fu_acc_0_31017_37376 : unsigned (7 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_335_i0_fu_acc_0_31017_37304 : unsigned (25 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_336_i0_fu_acc_0_31017_37313 : unsigned (24 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_337_i0_fu_acc_0_31017_37398 : unsigned (7 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_337_i1_fu_acc_0_31017_37409 : unsigned (7 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_338_i0_fu_acc_0_31017_37905 : unsigned (9 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_338_i1_fu_acc_0_31017_37932 : unsigned (9 downto 0);
  signal out_ui_rshift_expr_FU_32_0_32_339_i0_fu_acc_0_31017_37929 : unsigned (9 downto 0);
  signal out_ui_rshift_expr_FU_64_0_64_340_i0_fu_acc_0_31017_37737 : unsigned (22 downto 0);
  signal out_ui_rshift_expr_FU_64_0_64_341_i0_fu_acc_0_31017_37752 : unsigned (22 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i0_fu_acc_0_31017_36874 : unsigned (5 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i1_fu_acc_0_31017_36922 : unsigned (6 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i2_fu_acc_0_31017_36925 : unsigned (6 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i3_fu_acc_0_31017_36928 : unsigned (5 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i4_fu_acc_0_31017_36931 : unsigned (5 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i5_fu_acc_0_31017_37075 : unsigned (1 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i6_fu_acc_0_31017_37096 : unsigned (2 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_342_i7_fu_acc_0_31017_37102 : unsigned (1 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_343_i0_fu_acc_0_31017_37060 : unsigned (5 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_344_i0_fu_acc_0_31017_37593 : unsigned (0 downto 0);
  signal out_ui_rshift_expr_FU_8_0_8_344_i1_fu_acc_0_31017_37662 : unsigned (0 downto 0);
  signal out_ui_ternary_plus_expr_FU_0_16_16_16_345_i0_fu_acc_0_31017_37611 : unsigned (9 downto 0);
  signal out_vb_assign_conn_obj_2_ASSIGN_VECTOR_BOOL_FU_vb_assign_2 : std_logic_vector(31 downto 0) ;
  signal s_MEMORY_CTRL_D21_251_i00 : std_logic;
  signal s_done_MEMORY_CTRL_D21_251_i0 : std_logic;
  signal sig_in_bus_mergerMout_Wdata_ram0_0 : std_logic_vector(31 downto 0) ;
  signal sig_in_bus_mergerMout_addr_ram1_0 : std_logic_vector(31 downto 0) ;
  signal sig_in_bus_mergerMout_data_ram_size2_0 : std_logic_vector(5 downto 0) ;
  signal sig_in_bus_mergerMout_oe_ram3_0 : std_logic;
  signal sig_in_bus_mergerMout_we_ram4_0 : std_logic;
  signal \sig_out_bus_mergerMout_Wdata_ram0_\ : std_logic_vector(31 downto 0) ;
  signal \sig_out_bus_mergerMout_addr_ram1_\ : std_logic_vector(31 downto 0) ;
  signal \sig_out_bus_mergerMout_data_ram_size2_\ : std_logic_vector(5 downto 0) ;
  signal \sig_out_bus_mergerMout_oe_ram3_\ : std_logic_vector(0 downto 0);
  signal \sig_out_bus_mergerMout_we_ram4_\ : std_logic_vector(0 downto 0);
begin
  ASSIGN_VECTOR_BOOL_FU_vb_assign_2 : ASSIGN_VECTOR_BOOL_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_vb_assign_conn_obj_2_ASSIGN_VECTOR_BOOL_FU_vb_assign_2,
    in1 => out_reg_47_reg_47);
  IUdata_converter_FU_iu_conv_0 : IUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_iu_conv_conn_obj_0_IUdata_converter_FU_iu_conv_0,
    in1 => signed(out_reg_18_reg_18));
  IUdata_converter_FU_iu_conv_1 : IUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_iu_conv_conn_obj_1_IUdata_converter_FU_iu_conv_1,
    in1 => signed(out_reg_17_reg_17));
  MEMORY_CTRL_D21_251_i0 : MEMORY_CTRL_D21 generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_in3=>6,
    BITSIZE_out1=>32,
    BITSIZE_Min_addr_ram=>32,
    BITSIZE_Mout_addr_ram=>32,
    BITSIZE_M_Rdata_ram=>32,
    BITSIZE_Min_Wdata_ram=>32,
    BITSIZE_Mout_Wdata_ram=>32,
    BITSIZE_Min_data_ram_size=>6,
    BITSIZE_Mout_data_ram_size=>6) port map (done_port => s_done_MEMORY_CTRL_D21_251_i0,
    out1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    Mout_oe_ram => sig_in_bus_mergerMout_oe_ram3_0,
    Mout_we_ram => sig_in_bus_mergerMout_we_ram4_0,
    Mout_addr_ram => sig_in_bus_mergerMout_addr_ram1_0,
    Mout_Wdata_ram => sig_in_bus_mergerMout_Wdata_ram0_0,
    Mout_data_ram_size => sig_in_bus_mergerMout_data_ram_size2_0,
    clock => clock,
    start_port => s_MEMORY_CTRL_D21_251_i00,
    in1 => out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1,
    in2 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0,
    in3 => out_conv_out_const_6_7_6,
    in4 => out_const_15(0),
    sel_LOAD => fuselector_MEMORY_CTRL_D21_251_i0_LOAD,
    sel_STORE => fuselector_MEMORY_CTRL_D21_251_i0_STORE,
    Min_oe_ram => Min_oe_ram,
    Min_we_ram => Min_we_ram,
    Min_addr_ram => Min_addr_ram,
    M_Rdata_ram => M_Rdata_ram,
    Min_Wdata_ram => Min_Wdata_ram,
    Min_data_ram_size => Min_data_ram_size,
    M_DataRdy => M_DataRdy);
  MUX_550_reg_13_0_0_0 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_550_reg_13_0_0_0,
    sel => selector_MUX_550_reg_13_0_0_0,
    in1 => std_logic_vector(out_ui_bit_ior_concat_expr_FU_277_i0_fu_acc_0_31017_37385),
    in2 => std_logic_vector(out_ui_lshift_expr_FU_32_0_32_296_i0_fu_acc_0_31017_36844));
  MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0,
    sel => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0,
    in1 => std_logic_vector(out_iu_conv_conn_obj_0_IUdata_converter_FU_iu_conv_0),
    in2 => std_logic_vector(out_iu_conv_conn_obj_1_IUdata_converter_FU_iu_conv_1));
  MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1,
    sel => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1,
    in1 => out_vb_assign_conn_obj_2_ASSIGN_VECTOR_BOOL_FU_vb_assign_2,
    in2 => out_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0,
    in1 => out_reg_8_reg_8,
    in2 => out_reg_7_reg_7);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1,
    in1 => out_reg_6_reg_6,
    in2 => out_reg_5_reg_5);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2,
    in1 => out_reg_4_reg_4,
    in2 => out_reg_3_reg_3);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3,
    in1 => out_reg_2_reg_2,
    in2 => out_reg_19_reg_19);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4,
    in1 => out_reg_1_reg_1,
    in2 => out_UUdata_converter_FU_3_i0_fu_acc_0_31017_31446);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0,
    in1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0,
    in2 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1,
    in1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2,
    in2 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2,
    in1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4,
    in2 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0);
  MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : MUX_GATE generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0,
    sel => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0,
    in1 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1,
    in2 => out_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2);
  \bus_mergerMout_Wdata_ram0_\ : bus_merger generic map(BITSIZE_in1=>32, PORTSIZE_in1=>1,
    BITSIZE_out1=>32) port map (out1 => \sig_out_bus_mergerMout_Wdata_ram0_\,
      in1(31 downto 0) => sig_in_bus_mergerMout_Wdata_ram0_0);
  \bus_mergerMout_addr_ram1_\ : bus_merger generic map(BITSIZE_in1=>32, PORTSIZE_in1=>1,
    BITSIZE_out1=>32) port map (out1 => \sig_out_bus_mergerMout_addr_ram1_\,
      in1(31 downto 0) => sig_in_bus_mergerMout_addr_ram1_0);
  \bus_mergerMout_data_ram_size2_\ : bus_merger generic map(BITSIZE_in1=>6, PORTSIZE_in1=>1,
    BITSIZE_out1=>6) port map (out1 => \sig_out_bus_mergerMout_data_ram_size2_\,
      in1(5 downto 0) => sig_in_bus_mergerMout_data_ram_size2_0);
  \bus_mergerMout_oe_ram3_\ : bus_merger generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => \sig_out_bus_mergerMout_oe_ram3_\,
      in1(0) => sig_in_bus_mergerMout_oe_ram3_0);
  \bus_mergerMout_we_ram4_\ : bus_merger generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => \sig_out_bus_mergerMout_we_ram4_\,
      in1(0) => sig_in_bus_mergerMout_we_ram4_0);
  const_0 : constant_value generic map(BITSIZE_out1=>1,
    value=>"0") port map (out1 => out_const_0);
  const_1 : constant_value generic map(BITSIZE_out1=>2,
    value=>"01") port map (out1 => out_const_1);
  const_10 : constant_value generic map(BITSIZE_out1=>5,
    value=>"01100") port map (out1 => out_const_10);
  const_11 : constant_value generic map(BITSIZE_out1=>6,
    value=>"011000") port map (out1 => out_const_11);
  const_12 : constant_value generic map(BITSIZE_out1=>6,
    value=>"011001") port map (out1 => out_const_12);
  const_13 : constant_value generic map(BITSIZE_out1=>4,
    value=>"0111") port map (out1 => out_const_13);
  const_14 : constant_value generic map(BITSIZE_out1=>6,
    value=>"011111") port map (out1 => out_const_14);
  const_15 : constant_value generic map(BITSIZE_out1=>1,
    value=>"1") port map (out1 => out_const_15);
  const_16 : constant_value generic map(BITSIZE_out1=>2,
    value=>"10") port map (out1 => out_const_16);
  const_17 : constant_value generic map(BITSIZE_out1=>3,
    value=>"100") port map (out1 => out_const_17);
  const_18 : constant_value generic map(BITSIZE_out1=>4,
    value=>"1000") port map (out1 => out_const_18);
  const_19 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10000") port map (out1 => out_const_19);
  const_2 : constant_value generic map(BITSIZE_out1=>3,
    value=>"010") port map (out1 => out_const_2);
  const_20 : constant_value generic map(BITSIZE_out1=>6,
    value=>"100000") port map (out1 => out_const_20);
  const_21 : constant_value generic map(BITSIZE_out1=>8,
    value=>"10000000") port map (out1 => out_const_21);
  const_22 : constant_value generic map(BITSIZE_out1=>17,
    value=>"10000000000000000") port map (out1 => out_const_22);
  const_23 : constant_value generic map(BITSIZE_out1=>24,
    value=>"100000000000000000000000") port map (out1 => out_const_23);
  const_24 : constant_value generic map(BITSIZE_out1=>32,
    value=>"10000000000000000000000000000000") port map (out1 => out_const_24);
  const_25 : constant_value generic map(BITSIZE_out1=>33,
    value=>"100000000000000000000000000000000") port map (out1 => out_const_25);
  const_26 : constant_value generic map(BITSIZE_out1=>64,
    value=>"1000000000000000000000000000000000000000000000000000000000000000") port map (out1 => out_const_26);
  const_27 : constant_value generic map(BITSIZE_out1=>49,
    value=>"1000000000000111100010001000100011111111111111111") port map (out1 => out_const_27);
  const_28 : constant_value generic map(BITSIZE_out1=>59,
    value=>"10000010101100011001001110100100110001101111010111010111111") port map (out1 => out_const_28);
  const_29 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10001") port map (out1 => out_const_29);
  const_3 : constant_value generic map(BITSIZE_out1=>4,
    value=>"0100") port map (out1 => out_const_3);
  const_30 : constant_value generic map(BITSIZE_out1=>61,
    value=>"1000100010001000000000000111100010001000100010000000000000000") port map (out1 => out_const_30);
  const_31 : constant_value generic map(BITSIZE_out1=>4,
    value=>"1001") port map (out1 => out_const_31);
  const_32 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10011") port map (out1 => out_const_32);
  const_33 : constant_value generic map(BITSIZE_out1=>3,
    value=>"101") port map (out1 => out_const_33);
  const_34 : constant_value generic map(BITSIZE_out1=>27,
    value=>"101000001010000000000110011") port map (out1 => out_const_34);
  const_35 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10101") port map (out1 => out_const_35);
  const_36 : constant_value generic map(BITSIZE_out1=>64,
    value=>"1010101010101010110011001100110011110000111100001111111100000000") port map (out1 => out_const_36);
  const_37 : constant_value generic map(BITSIZE_out1=>48,
    value=>"101011001111111100000000000000001010110000000000") port map (out1 => out_const_37);
  const_38 : constant_value generic map(BITSIZE_out1=>4,
    value=>"1011") port map (out1 => out_const_38);
  const_39 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10110") port map (out1 => out_const_39);
  const_4 : constant_value generic map(BITSIZE_out1=>5,
    value=>"01000") port map (out1 => out_const_4);
  const_40 : constant_value generic map(BITSIZE_out1=>5,
    value=>"10111") port map (out1 => out_const_40);
  const_41 : constant_value generic map(BITSIZE_out1=>6,
    value=>"101111") port map (out1 => out_const_41);
  const_42 : constant_value generic map(BITSIZE_out1=>2,
    value=>"11") port map (out1 => out_const_42);
  const_43 : constant_value generic map(BITSIZE_out1=>3,
    value=>"110") port map (out1 => out_const_43);
  const_44 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11000") port map (out1 => out_const_44);
  const_45 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11001") port map (out1 => out_const_45);
  const_46 : constant_value generic map(BITSIZE_out1=>8,
    value=>"11001111") port map (out1 => out_const_46);
  const_47 : constant_value generic map(BITSIZE_out1=>4,
    value=>"1101") port map (out1 => out_const_47);
  const_48 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11010") port map (out1 => out_const_48);
  const_49 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11011") port map (out1 => out_const_49);
  const_5 : constant_value generic map(BITSIZE_out1=>6,
    value=>"010000") port map (out1 => out_const_5);
  const_50 : constant_value generic map(BITSIZE_out1=>8,
    value=>"11011000") port map (out1 => out_const_50);
  const_51 : constant_value generic map(BITSIZE_out1=>3,
    value=>"111") port map (out1 => out_const_51);
  const_52 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11100") port map (out1 => out_const_52);
  const_53 : constant_value generic map(BITSIZE_out1=>8,
    value=>"11100000") port map (out1 => out_const_53);
  const_54 : constant_value generic map(BITSIZE_out1=>56,
    value=>"11100000000000000000000011111111000111111111111111111111") port map (out1 => out_const_54);
  const_55 : constant_value generic map(BITSIZE_out1=>12,
    value=>"111000001111") port map (out1 => out_const_55);
  const_56 : constant_value generic map(BITSIZE_out1=>11,
    value=>"11100001111") port map (out1 => out_const_56);
  const_57 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11101") port map (out1 => out_const_57);
  const_58 : constant_value generic map(BITSIZE_out1=>8,
    value=>"11101010") port map (out1 => out_const_58);
  const_59 : constant_value generic map(BITSIZE_out1=>4,
    value=>"1111") port map (out1 => out_const_59);
  const_6 : constant_value generic map(BITSIZE_out1=>7,
    value=>"0100000") port map (out1 => out_const_6);
  const_60 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11110") port map (out1 => out_const_60);
  const_61 : constant_value generic map(BITSIZE_out1=>32,
    value=>"11110111101000101101010110000000") port map (out1 => out_const_61);
  const_62 : constant_value generic map(BITSIZE_out1=>5,
    value=>"11111") port map (out1 => out_const_62);
  const_63 : constant_value generic map(BITSIZE_out1=>32,
    value=>"11111010111110101111111111001100") port map (out1 => out_const_63);
  const_64 : constant_value generic map(BITSIZE_out1=>6,
    value=>"111111") port map (out1 => out_const_64);
  const_65 : constant_value generic map(BITSIZE_out1=>8,
    value=>"11111111") port map (out1 => out_const_65);
  const_66 : constant_value generic map(BITSIZE_out1=>31,
    value=>"1111111100000000000000000000000") port map (out1 => out_const_66);
  const_67 : constant_value generic map(BITSIZE_out1=>10,
    value=>"1111111111") port map (out1 => out_const_67);
  const_68 : constant_value generic map(BITSIZE_out1=>48,
    value=>"111111111111111000000000000000000000000000000000") port map (out1 => out_const_68);
  const_69 : constant_value generic map(BITSIZE_out1=>64,
    value=>"1111111111111110000000000000000000000000000000000000000000000000") port map (out1 => out_const_69);
  const_7 : constant_value generic map(BITSIZE_out1=>9,
    value=>"010011100") port map (out1 => out_const_7);
  const_70 : constant_value generic map(BITSIZE_out1=>17,
    value=>"11111111111111110") port map (out1 => out_const_70);
  const_71 : constant_value generic map(BITSIZE_out1=>17,
    value=>"11111111111111111") port map (out1 => out_const_71);
  const_72 : constant_value generic map(BITSIZE_out1=>32,
    value=>"11111111111111111010110000000000") port map (out1 => out_const_72);
  const_73 : constant_value generic map(BITSIZE_out1=>23,
    value=>"11111111111111111111111") port map (out1 => out_const_73);
  const_74 : constant_value generic map(BITSIZE_out1=>32,
    value=>"11111111111111111111111110000001") port map (out1 => out_const_74);
  const_75 : constant_value generic map(BITSIZE_out1=>31,
    value=>"1111111111111111111111111111111") port map (out1 => out_const_75);
  const_76 : constant_value generic map(BITSIZE_out1=>32,
    value=>"11111111111111111111111111111111") port map (out1 => out_const_76);
  const_77 : constant_value generic map(BITSIZE_out1=>33,
    value=>"111111111111111111111111111111111") port map (out1 => out_const_77);
  const_78 : constant_value generic map(BITSIZE_out1=>47,
    value=>"11111111111111111111111111111111111111111111111") port map (out1 => out_const_78);
  const_8 : constant_value generic map(BITSIZE_out1=>6,
    value=>"010100") port map (out1 => out_const_8);
  const_9 : constant_value generic map(BITSIZE_out1=>6,
    value=>"010111") port map (out1 => out_const_9);
  conv_out_const_6_7_6 : UUdata_converter_FU generic map(BITSIZE_in1=>7,
    BITSIZE_out1=>6) port map (out1 => out_conv_out_const_6_7_6,
    in1 => out_const_6);
  fu_acc_0_31017_31058 : plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_plus_expr_FU_32_32_32_260_i0_fu_acc_0_31017_31058,
    in1 => signed(out_reg_0_reg_0),
    in2 => signed(out_reg_9_reg_9));
  fu_acc_0_31017_31062 : mult_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32,
    PIPE_PARAMETER=>0) port map (out1 => out_mult_expr_FU_32_32_32_0_258_i0_fu_acc_0_31017_31062,
    clock => clock,
    in1 => signed(out_reg_9_reg_9),
    in2 => signed(out_reg_10_reg_10));
  fu_acc_0_31017_31446 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_3_i0_fu_acc_0_31017_31446,
    in1 => out_UUdata_converter_FU_2_i0_fu_acc_0_31017_31544);
  fu_acc_0_31017_31466 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_5_i0_fu_acc_0_31017_31466,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_321_i0_fu_acc_0_31017_31564));
  fu_acc_0_31017_31479 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_7_i0_fu_acc_0_31017_31479,
    in1 => out_UUdata_converter_FU_6_i0_fu_acc_0_31017_31573);
  fu_acc_0_31017_31492 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_9_i0_fu_acc_0_31017_31492,
    in1 => out_UUdata_converter_FU_8_i0_fu_acc_0_31017_31585);
  fu_acc_0_31017_31501 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_320_i0_fu_acc_0_31017_31501,
    in1 => unsigned(out_UUdata_converter_FU_9_i0_fu_acc_0_31017_31492),
    in2 => unsigned(out_const_17));
  fu_acc_0_31017_31505 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_11_i0_fu_acc_0_31017_31505,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_321_i1_fu_acc_0_31017_31600));
  fu_acc_0_31017_31514 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_320_i1_fu_acc_0_31017_31514,
    in1 => unsigned(out_UUdata_converter_FU_11_i0_fu_acc_0_31017_31505),
    in2 => unsigned(out_const_17));
  fu_acc_0_31017_31518 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_13_i0_fu_acc_0_31017_31518,
    in1 => out_UUdata_converter_FU_12_i0_fu_acc_0_31017_31609);
  fu_acc_0_31017_31527 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_320_i2_fu_acc_0_31017_31527,
    in1 => unsigned(out_UUdata_converter_FU_13_i0_fu_acc_0_31017_31518),
    in2 => unsigned(out_const_17));
  fu_acc_0_31017_31544 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_2_i0_fu_acc_0_31017_31544,
    in1 => in_port_param);
  fu_acc_0_31017_31560 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_4_i0_fu_acc_0_31017_31560,
    in1 => in_port_param);
  fu_acc_0_31017_31564 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_321_i0_fu_acc_0_31017_31564,
    in1 => unsigned(out_UUdata_converter_FU_4_i0_fu_acc_0_31017_31560),
    in2 => unsigned(out_const_18));
  fu_acc_0_31017_31573 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_6_i0_fu_acc_0_31017_31573,
    in1 => in_port_result);
  fu_acc_0_31017_31585 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_8_i0_fu_acc_0_31017_31585,
    in1 => in_port_param);
  fu_acc_0_31017_31597 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_10_i0_fu_acc_0_31017_31597,
    in1 => in_port_param);
  fu_acc_0_31017_31600 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_321_i1_fu_acc_0_31017_31600,
    in1 => unsigned(out_UUdata_converter_FU_10_i0_fu_acc_0_31017_31597),
    in2 => unsigned(out_const_18));
  fu_acc_0_31017_31609 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_12_i0_fu_acc_0_31017_31609,
    in1 => in_port_result);
  fu_acc_0_31017_31621 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_113_i0_fu_acc_0_31017_31621,
    in1 => in_port_param);
  fu_acc_0_31017_31625 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_322_i0_fu_acc_0_31017_31625,
    in1 => unsigned(out_UUdata_converter_FU_113_i0_fu_acc_0_31017_31621),
    in2 => unsigned(out_const_19));
  fu_acc_0_31017_31629 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_114_i0_fu_acc_0_31017_31629,
    in1 => in_port_result);
  fu_acc_0_31017_31632 : ui_pointer_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4,
    BITSIZE_out1=>32,
    LSB_PARAMETER=>0) port map (out1 => out_ui_pointer_plus_expr_FU_32_0_32_321_i2_fu_acc_0_31017_31632,
    in1 => unsigned(out_UUdata_converter_FU_114_i0_fu_acc_0_31017_31629),
    in2 => unsigned(out_const_18));
  fu_acc_0_31017_33175 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_238_i0_fu_acc_0_31017_33175,
    in1 => std_logic_vector(out_ui_cond_expr_FU_32_32_32_32_288_i6_fu_acc_0_31017_37941));
  fu_acc_0_31017_33178 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>31) port map (out1 => out_UUdata_converter_FU_117_i0_fu_acc_0_31017_33178,
    in1 => out_reg_13_reg_13);
  fu_acc_0_31017_33181 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>31) port map (out1 => out_UUdata_converter_FU_118_i0_fu_acc_0_31017_33181,
    in1 => out_reg_29_reg_29);
  fu_acc_0_31017_36800 : eq_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_eq_expr_FU_32_0_32_255_i0_fu_acc_0_31017_36800,
    in1 => signed(out_reg_9_reg_9),
    in2 => signed(out_const_0));
  fu_acc_0_31017_36805 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_14_i0_fu_acc_0_31017_36805,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_62);
  fu_acc_0_31017_36808 : eq_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>32,
    BITSIZE_out1=>1) port map (out1 => out_eq_expr_FU_32_0_32_256_i0_fu_acc_0_31017_36808,
    in1 => signed(out_reg_9_reg_9),
    in2 => signed(out_const_24));
  fu_acc_0_31017_36811 : IUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_15_i0_fu_acc_0_31017_36811,
    in1 => signed(out_reg_9_reg_9));
  fu_acc_0_31017_36814 : negate_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in1 => signed(out_reg_9_reg_9));
  fu_acc_0_31017_36817 : IUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_16_i0_fu_acc_0_31017_36817,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814);
  fu_acc_0_31017_36820 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_17_i0_fu_acc_0_31017_36820,
    in1(0) => out_extract_bit_expr_FU_14_i0_fu_acc_0_31017_36805);
  fu_acc_0_31017_36823 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>6,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_294_i0_fu_acc_0_31017_36823,
    in1 => unsigned(out_UUdata_converter_FU_17_i0_fu_acc_0_31017_36820),
    in2 => out_const_14);
  fu_acc_0_31017_36826 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>1,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_324_i0_fu_acc_0_31017_36826,
    in1 => out_ui_lshift_expr_FU_32_0_32_294_i0_fu_acc_0_31017_36823,
    in2 => out_const_62);
  fu_acc_0_31017_36829 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_295_i0_fu_acc_0_31017_36829,
    in1 => out_ui_rshift_expr_FU_32_0_32_324_i0_fu_acc_0_31017_36826,
    in2 => out_const_62);
  fu_acc_0_31017_36832 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_18_i0_fu_acc_0_31017_36832,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_62);
  fu_acc_0_31017_36835 : lut_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835,
    in1 => out_const_16,
    in2 => out_extract_bit_expr_FU_18_i0_fu_acc_0_31017_36832,
    in3 => out_eq_expr_FU_32_0_32_256_i0_fu_acc_0_31017_36808(0),
    in4 => out_eq_expr_FU_32_0_32_255_i0_fu_acc_0_31017_36800(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36838 : lut_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_20_i0_fu_acc_0_31017_36838,
    in1 => out_const_15,
    in2 => out_eq_expr_FU_32_0_32_256_i0_fu_acc_0_31017_36808(0),
    in3 => out_eq_expr_FU_32_0_32_255_i0_fu_acc_0_31017_36800(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36841 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_in3=>8,
    BITSIZE_out1=>8) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i0_fu_acc_0_31017_36841,
    in1 => out_eq_expr_FU_32_0_32_255_i0_fu_acc_0_31017_36800,
    in2 => unsigned(out_const_0),
    in3 => unsigned(out_const_46));
  fu_acc_0_31017_36844 : ui_lshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_296_i0_fu_acc_0_31017_36844,
    in1 => out_ui_cond_expr_FU_8_8_8_8_289_i0_fu_acc_0_31017_36841,
    in2 => out_const_44);
  fu_acc_0_31017_36847 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>32,
    BITSIZE_in3=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i0_fu_acc_0_31017_36847,
    in1 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835,
    in2 => out_IUdata_converter_FU_16_i0_fu_acc_0_31017_36817,
    in3 => out_IUdata_converter_FU_15_i0_fu_acc_0_31017_36811);
  fu_acc_0_31017_36850 : UUdata_converter_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850,
    in1 => std_logic_vector(out_ui_cond_expr_FU_32_32_32_32_288_i0_fu_acc_0_31017_36847));
  fu_acc_0_31017_36853 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>6,
    BITSIZE_out1=>16,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_325_i0_fu_acc_0_31017_36853,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_5);
  fu_acc_0_31017_36856 : ui_eq_expr_FU generic map(BITSIZE_in1=>16,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_16_0_16_290_i0_fu_acc_0_31017_36856,
    in1 => out_ui_rshift_expr_FU_32_0_32_325_i0_fu_acc_0_31017_36853,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36859 : ui_eq_expr_FU generic map(BITSIZE_in1=>16,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859,
    in1 => out_ui_rshift_expr_FU_32_0_32_325_i0_fu_acc_0_31017_36853,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36862 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>6,
    BITSIZE_out1=>8,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_326_i0_fu_acc_0_31017_36862,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_11);
  fu_acc_0_31017_36865 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>6,
    BITSIZE_out1=>12,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_327_i0_fu_acc_0_31017_36865,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_8);
  fu_acc_0_31017_36868 : ui_eq_expr_FU generic map(BITSIZE_in1=>12,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_16_0_16_290_i2_fu_acc_0_31017_36868,
    in1 => out_ui_rshift_expr_FU_32_0_32_327_i0_fu_acc_0_31017_36865,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36871 : ui_rshift_expr_FU generic map(BITSIZE_in1=>16,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_16_0_16_323_i0_fu_acc_0_31017_36871,
    in1 => out_ui_rshift_expr_FU_32_0_32_325_i0_fu_acc_0_31017_36853,
    in2 => out_const_15);
  fu_acc_0_31017_36874 : ui_rshift_expr_FU generic map(BITSIZE_in1=>7,
    BITSIZE_in2=>1,
    BITSIZE_out1=>6,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i0_fu_acc_0_31017_36874,
    in1 => out_ui_rshift_expr_FU_16_0_16_323_i0_fu_acc_0_31017_36871,
    in2 => out_const_15);
  fu_acc_0_31017_36877 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>6,
    BITSIZE_in2=>6,
    BITSIZE_out1=>6) port map (out1 => out_ui_bit_and_expr_FU_8_0_8_272_i0_fu_acc_0_31017_36877,
    in1 => out_ui_rshift_expr_FU_8_0_8_342_i0_fu_acc_0_31017_36874,
    in2 => unsigned(out_const_64));
  fu_acc_0_31017_36880 : ui_lshift_expr_FU generic map(BITSIZE_in1=>6,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i0_fu_acc_0_31017_36880,
    in1 => out_ui_bit_and_expr_FU_8_0_8_272_i0_fu_acc_0_31017_36877,
    in2 => out_const_15);
  fu_acc_0_31017_36883 : ui_lshift_expr_FU generic map(BITSIZE_in1=>7,
    BITSIZE_in2=>1,
    BITSIZE_out1=>8,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i1_fu_acc_0_31017_36883,
    in1 => out_ui_lshift_expr_FU_8_0_8_307_i0_fu_acc_0_31017_36880,
    in2 => out_const_15);
  fu_acc_0_31017_36886 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>24,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_328_i0_fu_acc_0_31017_36886,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_4);
  fu_acc_0_31017_36889 : ui_eq_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889,
    in1 => out_ui_rshift_expr_FU_32_0_32_328_i0_fu_acc_0_31017_36886,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36892 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>20,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_329_i0_fu_acc_0_31017_36892,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_10);
  fu_acc_0_31017_36895 : ui_eq_expr_FU generic map(BITSIZE_in1=>20,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i1_fu_acc_0_31017_36895,
    in1 => out_ui_rshift_expr_FU_32_0_32_329_i0_fu_acc_0_31017_36892,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36898 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4,
    BITSIZE_out1=>28,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_330_i0_fu_acc_0_31017_36898,
    in1 => unsigned(out_UUdata_converter_FU_21_i0_fu_acc_0_31017_36850),
    in2 => out_const_3);
  fu_acc_0_31017_36901 : ui_eq_expr_FU generic map(BITSIZE_in1=>28,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i2_fu_acc_0_31017_36901,
    in1 => out_ui_rshift_expr_FU_32_0_32_330_i0_fu_acc_0_31017_36898,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_36904 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>8,
    BITSIZE_out1=>8) port map (out1 => out_ui_bit_and_expr_FU_8_0_8_273_i0_fu_acc_0_31017_36904,
    in1 => out_ui_cond_expr_FU_32_32_32_32_288_i0_fu_acc_0_31017_36847,
    in2 => unsigned(out_const_65));
  fu_acc_0_31017_36907 : UUdata_converter_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>8) port map (out1 => out_UUdata_converter_FU_22_i0_fu_acc_0_31017_36907,
    in1 => std_logic_vector(out_ui_bit_and_expr_FU_8_0_8_273_i0_fu_acc_0_31017_36904));
  fu_acc_0_31017_36910 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_23_i0_fu_acc_0_31017_36910,
    in1 => out_ui_eq_expr_FU_16_0_16_290_i0_fu_acc_0_31017_36856);
  fu_acc_0_31017_36913 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>4,
    BITSIZE_out1=>5,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_308_i0_fu_acc_0_31017_36913,
    in1 => unsigned(out_UUdata_converter_FU_23_i0_fu_acc_0_31017_36910),
    in2 => out_const_3);
  fu_acc_0_31017_36916 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916,
    in1 => out_const_18,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36919 : lut_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919,
    in1 => out_const_16,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36922 : ui_rshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i1_fu_acc_0_31017_36922,
    in1 => unsigned(out_UUdata_converter_FU_22_i0_fu_acc_0_31017_36907),
    in2 => out_const_15);
  fu_acc_0_31017_36925 : ui_rshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i2_fu_acc_0_31017_36925,
    in1 => out_ui_lshift_expr_FU_8_0_8_307_i1_fu_acc_0_31017_36883,
    in2 => out_const_15);
  fu_acc_0_31017_36928 : ui_rshift_expr_FU generic map(BITSIZE_in1=>7,
    BITSIZE_in2=>1,
    BITSIZE_out1=>6,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i3_fu_acc_0_31017_36928,
    in1 => out_ui_rshift_expr_FU_8_0_8_342_i1_fu_acc_0_31017_36922,
    in2 => out_const_15);
  fu_acc_0_31017_36931 : ui_rshift_expr_FU generic map(BITSIZE_in1=>7,
    BITSIZE_in2=>1,
    BITSIZE_out1=>6,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i4_fu_acc_0_31017_36931,
    in1 => out_ui_rshift_expr_FU_8_0_8_342_i2_fu_acc_0_31017_36925,
    in2 => out_const_15);
  fu_acc_0_31017_36934 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>6,
    BITSIZE_in3=>6,
    BITSIZE_out1=>6) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i1_fu_acc_0_31017_36934,
    in1 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916,
    in2 => out_ui_rshift_expr_FU_8_0_8_342_i3_fu_acc_0_31017_36928,
    in3 => out_ui_rshift_expr_FU_8_0_8_342_i4_fu_acc_0_31017_36931);
  fu_acc_0_31017_36937 : ui_lshift_expr_FU generic map(BITSIZE_in1=>6,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i2_fu_acc_0_31017_36937,
    in1 => out_ui_cond_expr_FU_8_8_8_8_289_i1_fu_acc_0_31017_36934,
    in2 => out_const_15);
  fu_acc_0_31017_36940 : ui_lshift_expr_FU generic map(BITSIZE_in1=>7,
    BITSIZE_in2=>1,
    BITSIZE_out1=>8,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i3_fu_acc_0_31017_36940,
    in1 => out_ui_lshift_expr_FU_8_0_8_307_i2_fu_acc_0_31017_36937,
    in2 => out_const_15);
  fu_acc_0_31017_36943 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_26_i0_fu_acc_0_31017_36943,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_44);
  fu_acc_0_31017_36946 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_27_i0_fu_acc_0_31017_36946,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_44);
  fu_acc_0_31017_36949 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_28_i0_fu_acc_0_31017_36949,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_45);
  fu_acc_0_31017_36952 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_29_i0_fu_acc_0_31017_36952,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_45);
  fu_acc_0_31017_36955 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_30_i0_fu_acc_0_31017_36955,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_48);
  fu_acc_0_31017_36958 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_31_i0_fu_acc_0_31017_36958,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_48);
  fu_acc_0_31017_36961 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_32_i0_fu_acc_0_31017_36961,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_49);
  fu_acc_0_31017_36964 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_33_i0_fu_acc_0_31017_36964,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_49);
  fu_acc_0_31017_36967 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_34_i0_fu_acc_0_31017_36967,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_52);
  fu_acc_0_31017_36970 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_35_i0_fu_acc_0_31017_36970,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_52);
  fu_acc_0_31017_36973 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_36_i0_fu_acc_0_31017_36973,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_57);
  fu_acc_0_31017_36976 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_37_i0_fu_acc_0_31017_36976,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_57);
  fu_acc_0_31017_36979 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_38_i0_fu_acc_0_31017_36979,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_60);
  fu_acc_0_31017_36982 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_39_i0_fu_acc_0_31017_36982,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_60);
  fu_acc_0_31017_36985 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_40_i0_fu_acc_0_31017_36985,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_62);
  fu_acc_0_31017_36988 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_41_i0_fu_acc_0_31017_36988,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_62);
  fu_acc_0_31017_36991 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_42_i0_fu_acc_0_31017_36991,
    in1 => out_const_63,
    in2 => out_extract_bit_expr_FU_30_i0_fu_acc_0_31017_36955,
    in3 => out_extract_bit_expr_FU_31_i0_fu_acc_0_31017_36958,
    in4 => out_extract_bit_expr_FU_32_i0_fu_acc_0_31017_36961,
    in5 => out_extract_bit_expr_FU_33_i0_fu_acc_0_31017_36964,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36994 : lut_expr_FU generic map(BITSIZE_in1=>27,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_43_i0_fu_acc_0_31017_36994,
    in1 => out_const_34,
    in2 => out_extract_bit_expr_FU_26_i0_fu_acc_0_31017_36943,
    in3 => out_extract_bit_expr_FU_27_i0_fu_acc_0_31017_36946,
    in4 => out_extract_bit_expr_FU_28_i0_fu_acc_0_31017_36949,
    in5 => out_extract_bit_expr_FU_29_i0_fu_acc_0_31017_36952,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_42_i0_fu_acc_0_31017_36991(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_36997 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_44_i0_fu_acc_0_31017_36997,
    in1 => out_const_63,
    in2 => out_extract_bit_expr_FU_38_i0_fu_acc_0_31017_36979,
    in3 => out_extract_bit_expr_FU_39_i0_fu_acc_0_31017_36982,
    in4 => out_extract_bit_expr_FU_40_i0_fu_acc_0_31017_36985,
    in5 => out_extract_bit_expr_FU_41_i0_fu_acc_0_31017_36988,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37000 : lut_expr_FU generic map(BITSIZE_in1=>27,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_45_i0_fu_acc_0_31017_37000,
    in1 => out_const_34,
    in2 => out_extract_bit_expr_FU_34_i0_fu_acc_0_31017_36967,
    in3 => out_extract_bit_expr_FU_35_i0_fu_acc_0_31017_36970,
    in4 => out_extract_bit_expr_FU_36_i0_fu_acc_0_31017_36973,
    in5 => out_extract_bit_expr_FU_37_i0_fu_acc_0_31017_36976,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_44_i0_fu_acc_0_31017_36997(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37003 : lut_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_46_i0_fu_acc_0_31017_37003,
    in1 => out_const_58,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_lut_expr_FU_43_i0_fu_acc_0_31017_36994(0),
    in4 => out_lut_expr_FU_45_i0_fu_acc_0_31017_37000(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37006 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>24,
    BITSIZE_in3=>8,
    BITSIZE_out1=>24) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i1_fu_acc_0_31017_37006,
    in1 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919,
    in2 => out_ui_rshift_expr_FU_32_0_32_328_i0_fu_acc_0_31017_36886,
    in3 => out_ui_lshift_expr_FU_8_0_8_307_i3_fu_acc_0_31017_36940);
  fu_acc_0_31017_37009 : lut_expr_FU generic map(BITSIZE_in1=>5,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009,
    in1 => out_const_35,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_lut_expr_FU_43_i0_fu_acc_0_31017_36994(0),
    in4 => out_lut_expr_FU_45_i0_fu_acc_0_31017_37000(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37012 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_48_i0_fu_acc_0_31017_37012,
    in1 => out_const_47,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889(0),
    in4 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37015 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_49_i0_fu_acc_0_31017_37015,
    in1 => out_lut_expr_FU_48_i0_fu_acc_0_31017_37012);
  fu_acc_0_31017_37018 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_out1=>4,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_309_i0_fu_acc_0_31017_37018,
    in1 => unsigned(out_UUdata_converter_FU_49_i0_fu_acc_0_31017_37015),
    in2 => out_const_42);
  fu_acc_0_31017_37021 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_50_i0_fu_acc_0_31017_37021,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_52);
  fu_acc_0_31017_37024 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_51_i0_fu_acc_0_31017_37024,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_52);
  fu_acc_0_31017_37027 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_52_i0_fu_acc_0_31017_37027,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_57);
  fu_acc_0_31017_37030 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_53_i0_fu_acc_0_31017_37030,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_57);
  fu_acc_0_31017_37033 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_54_i0_fu_acc_0_31017_37033,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_60);
  fu_acc_0_31017_37036 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_55_i0_fu_acc_0_31017_37036,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_60);
  fu_acc_0_31017_37039 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_56_i0_fu_acc_0_31017_37039,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_62);
  fu_acc_0_31017_37042 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_57_i0_fu_acc_0_31017_37042,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_62);
  fu_acc_0_31017_37045 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_58_i0_fu_acc_0_31017_37045,
    in1 => out_const_63,
    in2 => out_extract_bit_expr_FU_50_i0_fu_acc_0_31017_37021,
    in3 => out_extract_bit_expr_FU_51_i0_fu_acc_0_31017_37024,
    in4 => out_extract_bit_expr_FU_52_i0_fu_acc_0_31017_37027,
    in5 => out_extract_bit_expr_FU_53_i0_fu_acc_0_31017_37030,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37048 : lut_expr_FU generic map(BITSIZE_in1=>27,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_59_i0_fu_acc_0_31017_37048,
    in1 => out_const_34,
    in2 => out_extract_bit_expr_FU_54_i0_fu_acc_0_31017_37033,
    in3 => out_extract_bit_expr_FU_55_i0_fu_acc_0_31017_37036,
    in4 => out_extract_bit_expr_FU_56_i0_fu_acc_0_31017_37039,
    in5 => out_extract_bit_expr_FU_57_i0_fu_acc_0_31017_37042,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_58_i0_fu_acc_0_31017_37045(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37051 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_60_i0_fu_acc_0_31017_37051,
    in1 => out_const_61,
    in2 => out_ui_eq_expr_FU_16_0_16_290_i1_fu_acc_0_31017_36859(0),
    in3 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_acc_0_31017_36889(0),
    in4 => out_ui_eq_expr_FU_32_0_32_291_i2_fu_acc_0_31017_36901(0),
    in5 => out_ui_eq_expr_FU_16_0_16_290_i2_fu_acc_0_31017_36868(0),
    in6 => out_ui_eq_expr_FU_32_0_32_291_i1_fu_acc_0_31017_36895(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37054 : lut_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_61_i0_fu_acc_0_31017_37054,
    in1 => out_const_50,
    in2 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in3 => out_lut_expr_FU_59_i0_fu_acc_0_31017_37048(0),
    in4 => out_lut_expr_FU_60_i0_fu_acc_0_31017_37051(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37057 : ui_rshift_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>2,
    BITSIZE_out1=>22,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_331_i0_fu_acc_0_31017_37057,
    in1 => out_ui_cond_expr_FU_32_32_32_32_288_i1_fu_acc_0_31017_37006,
    in2 => out_const_16);
  fu_acc_0_31017_37060 : ui_rshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>2,
    BITSIZE_out1=>6,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_343_i0_fu_acc_0_31017_37060,
    in1 => out_ui_rshift_expr_FU_32_0_32_326_i0_fu_acc_0_31017_36862,
    in2 => out_const_16);
  fu_acc_0_31017_37063 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>22,
    BITSIZE_in3=>6,
    BITSIZE_out1=>22) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i2_fu_acc_0_31017_37063,
    in1 => out_lut_expr_FU_46_i0_fu_acc_0_31017_37003,
    in2 => out_ui_rshift_expr_FU_32_0_32_331_i0_fu_acc_0_31017_37057,
    in3 => out_ui_rshift_expr_FU_8_0_8_343_i0_fu_acc_0_31017_37060);
  fu_acc_0_31017_37066 : ui_lshift_expr_FU generic map(BITSIZE_in1=>22,
    BITSIZE_in2=>2,
    BITSIZE_out1=>24,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_297_i0_fu_acc_0_31017_37066,
    in1 => out_ui_cond_expr_FU_32_32_32_32_288_i2_fu_acc_0_31017_37063,
    in2 => out_const_16);
  fu_acc_0_31017_37069 : ui_rshift_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>4,
    BITSIZE_out1=>20,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_330_i1_fu_acc_0_31017_37069,
    in1 => out_ui_lshift_expr_FU_32_0_32_297_i0_fu_acc_0_31017_37066,
    in2 => out_const_3);
  fu_acc_0_31017_37072 : ui_rshift_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>1,
    BITSIZE_out1=>3,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_332_i0_fu_acc_0_31017_37072,
    in1 => out_ui_lshift_expr_FU_32_0_32_297_i0_fu_acc_0_31017_37066,
    in2 => out_const_15);
  fu_acc_0_31017_37075 : ui_rshift_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_in2=>1,
    BITSIZE_out1=>2,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i5_fu_acc_0_31017_37075,
    in1 => out_ui_rshift_expr_FU_32_0_32_332_i0_fu_acc_0_31017_37072,
    in2 => out_const_15);
  fu_acc_0_31017_37078 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_bit_and_expr_FU_8_0_8_274_i0_fu_acc_0_31017_37078,
    in1 => out_ui_rshift_expr_FU_8_0_8_342_i5_fu_acc_0_31017_37075,
    in2 => unsigned(out_const_42));
  fu_acc_0_31017_37081 : ui_lshift_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1,
    BITSIZE_out1=>3,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i4_fu_acc_0_31017_37081,
    in1 => out_ui_bit_and_expr_FU_8_0_8_274_i0_fu_acc_0_31017_37078,
    in2 => out_const_15);
  fu_acc_0_31017_37084 : ui_lshift_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_in2=>1,
    BITSIZE_out1=>4,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_307_i5_fu_acc_0_31017_37084,
    in1 => out_ui_lshift_expr_FU_8_0_8_307_i4_fu_acc_0_31017_37081,
    in2 => out_const_15);
  fu_acc_0_31017_37087 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_62_i0_fu_acc_0_31017_37087,
    in1 => out_lut_expr_FU_61_i0_fu_acc_0_31017_37054);
  fu_acc_0_31017_37090 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>3,
    BITSIZE_out1=>3,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_310_i0_fu_acc_0_31017_37090,
    in1 => unsigned(out_UUdata_converter_FU_62_i0_fu_acc_0_31017_37087),
    in2 => out_const_2);
  fu_acc_0_31017_37093 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>5,
    BITSIZE_in2=>4,
    BITSIZE_out1=>5) port map (out1 => out_ui_bit_ior_expr_FU_0_8_8_282_i0_fu_acc_0_31017_37093,
    in1 => out_ui_lshift_expr_FU_8_0_8_308_i0_fu_acc_0_31017_36913,
    in2 => out_ui_lshift_expr_FU_8_0_8_309_i0_fu_acc_0_31017_37018);
  fu_acc_0_31017_37096 : ui_rshift_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_in2=>1,
    BITSIZE_out1=>3,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i6_fu_acc_0_31017_37096,
    in1 => out_ui_lshift_expr_FU_8_0_8_307_i5_fu_acc_0_31017_37084,
    in2 => out_const_15);
  fu_acc_0_31017_37099 : ui_rshift_expr_FU generic map(BITSIZE_in1=>20,
    BITSIZE_in2=>1,
    BITSIZE_out1=>19,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_332_i1_fu_acc_0_31017_37099,
    in1 => out_ui_rshift_expr_FU_32_0_32_330_i1_fu_acc_0_31017_37069,
    in2 => out_const_15);
  fu_acc_0_31017_37102 : ui_rshift_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_in2=>1,
    BITSIZE_out1=>2,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_8_0_8_342_i7_fu_acc_0_31017_37102,
    in1 => out_ui_rshift_expr_FU_8_0_8_342_i6_fu_acc_0_31017_37096,
    in2 => out_const_15);
  fu_acc_0_31017_37105 : ui_rshift_expr_FU generic map(BITSIZE_in1=>19,
    BITSIZE_in2=>1,
    BITSIZE_out1=>18,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_332_i2_fu_acc_0_31017_37105,
    in1 => out_ui_rshift_expr_FU_32_0_32_332_i1_fu_acc_0_31017_37099,
    in2 => out_const_15);
  fu_acc_0_31017_37108 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_in3=>18,
    BITSIZE_out1=>18) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i3_fu_acc_0_31017_37108,
    in1 => out_lut_expr_FU_61_i0_fu_acc_0_31017_37054,
    in2 => out_ui_rshift_expr_FU_8_0_8_342_i7_fu_acc_0_31017_37102,
    in3 => out_ui_rshift_expr_FU_32_0_32_332_i2_fu_acc_0_31017_37105);
  fu_acc_0_31017_37111 : ui_lshift_expr_FU generic map(BITSIZE_in1=>18,
    BITSIZE_in2=>1,
    BITSIZE_out1=>19,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_298_i0_fu_acc_0_31017_37111,
    in1 => out_ui_cond_expr_FU_32_32_32_32_288_i3_fu_acc_0_31017_37108,
    in2 => out_const_15);
  fu_acc_0_31017_37114 : ui_lshift_expr_FU generic map(BITSIZE_in1=>19,
    BITSIZE_in2=>1,
    BITSIZE_out1=>20,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_298_i1_fu_acc_0_31017_37114,
    in1 => out_ui_lshift_expr_FU_32_0_32_298_i0_fu_acc_0_31017_37111,
    in2 => out_const_15);
  fu_acc_0_31017_37117 : ui_rshift_expr_FU generic map(BITSIZE_in1=>20,
    BITSIZE_in2=>3,
    BITSIZE_out1=>18,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_333_i0_fu_acc_0_31017_37117,
    in1 => out_ui_lshift_expr_FU_32_0_32_298_i1_fu_acc_0_31017_37114,
    in2 => out_const_2);
  fu_acc_0_31017_37120 : ui_eq_expr_FU generic map(BITSIZE_in1=>18,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i3_fu_acc_0_31017_37120,
    in1 => out_ui_rshift_expr_FU_32_0_32_333_i0_fu_acc_0_31017_37117,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37123 : ui_eq_expr_FU generic map(BITSIZE_in1=>18,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i4_fu_acc_0_31017_37123,
    in1 => out_ui_rshift_expr_FU_32_0_32_333_i0_fu_acc_0_31017_37117,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37126 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_63_i0_fu_acc_0_31017_37126,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_38);
  fu_acc_0_31017_37129 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_64_i0_fu_acc_0_31017_37129,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_38);
  fu_acc_0_31017_37132 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>2) port map (out1 => out_extract_bit_expr_FU_65_i0_fu_acc_0_31017_37132,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_42);
  fu_acc_0_31017_37135 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>2) port map (out1 => out_extract_bit_expr_FU_66_i0_fu_acc_0_31017_37135,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_42);
  fu_acc_0_31017_37138 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_67_i0_fu_acc_0_31017_37138,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_32);
  fu_acc_0_31017_37141 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_68_i0_fu_acc_0_31017_37141,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_32);
  fu_acc_0_31017_37144 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_69_i0_fu_acc_0_31017_37144,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_49);
  fu_acc_0_31017_37147 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_70_i0_fu_acc_0_31017_37147,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_49);
  fu_acc_0_31017_37150 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_71_i0_fu_acc_0_31017_37150,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_59);
  fu_acc_0_31017_37153 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_72_i0_fu_acc_0_31017_37153,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_59);
  fu_acc_0_31017_37156 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_extract_bit_expr_FU_73_i0_fu_acc_0_31017_37156,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_51);
  fu_acc_0_31017_37159 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_extract_bit_expr_FU_74_i0_fu_acc_0_31017_37159,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_51);
  fu_acc_0_31017_37162 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_75_i0_fu_acc_0_31017_37162,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_40);
  fu_acc_0_31017_37165 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_76_i0_fu_acc_0_31017_37165,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_40);
  fu_acc_0_31017_37168 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_77_i0_fu_acc_0_31017_37168,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_62);
  fu_acc_0_31017_37171 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_78_i0_fu_acc_0_31017_37171,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_62);
  fu_acc_0_31017_37174 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_79_i0_fu_acc_0_31017_37174,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_31);
  fu_acc_0_31017_37177 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_80_i0_fu_acc_0_31017_37177,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_31);
  fu_acc_0_31017_37180 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_81_i0_fu_acc_0_31017_37180,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_15);
  fu_acc_0_31017_37183 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_82_i0_fu_acc_0_31017_37183,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_15);
  fu_acc_0_31017_37186 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_83_i0_fu_acc_0_31017_37186,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_29);
  fu_acc_0_31017_37189 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_84_i0_fu_acc_0_31017_37189,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_29);
  fu_acc_0_31017_37192 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_85_i0_fu_acc_0_31017_37192,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_45);
  fu_acc_0_31017_37195 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_86_i0_fu_acc_0_31017_37195,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_45);
  fu_acc_0_31017_37198 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_87_i0_fu_acc_0_31017_37198,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_47);
  fu_acc_0_31017_37201 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4) port map (out1 => out_extract_bit_expr_FU_88_i0_fu_acc_0_31017_37201,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_47);
  fu_acc_0_31017_37204 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_extract_bit_expr_FU_89_i0_fu_acc_0_31017_37204,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_33);
  fu_acc_0_31017_37207 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_extract_bit_expr_FU_90_i0_fu_acc_0_31017_37207,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_33);
  fu_acc_0_31017_37210 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_91_i0_fu_acc_0_31017_37210,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_35);
  fu_acc_0_31017_37213 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_92_i0_fu_acc_0_31017_37213,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_35);
  fu_acc_0_31017_37216 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_93_i0_fu_acc_0_31017_37216,
    in1 => out_negate_expr_FU_32_32_259_i0_fu_acc_0_31017_36814,
    in2 => out_const_57);
  fu_acc_0_31017_37219 : extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_extract_bit_expr_FU_94_i0_fu_acc_0_31017_37219,
    in1 => signed(out_reg_9_reg_9),
    in2 => out_const_57);
  fu_acc_0_31017_37222 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_95_i0_fu_acc_0_31017_37222,
    in1 => out_ui_eq_expr_FU_32_0_32_291_i3_fu_acc_0_31017_37120);
  fu_acc_0_31017_37225 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_8_0_8_311_i0_fu_acc_0_31017_37225,
    in1 => unsigned(out_UUdata_converter_FU_95_i0_fu_acc_0_31017_37222),
    in2 => out_const_1);
  fu_acc_0_31017_37228 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>3,
    BITSIZE_out1=>3) port map (out1 => out_ui_bit_ior_expr_FU_0_8_8_283_i0_fu_acc_0_31017_37228,
    in1 => out_ui_lshift_expr_FU_8_0_8_311_i0_fu_acc_0_31017_37225,
    in2 => out_ui_lshift_expr_FU_8_0_8_310_i0_fu_acc_0_31017_37090);
  fu_acc_0_31017_37231 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>5,
    BITSIZE_in2=>3,
    BITSIZE_out1=>5) port map (out1 => out_ui_bit_ior_expr_FU_0_8_8_284_i0_fu_acc_0_31017_37231,
    in1 => out_ui_bit_ior_expr_FU_0_8_8_282_i0_fu_acc_0_31017_37093,
    in2 => out_ui_bit_ior_expr_FU_0_8_8_283_i0_fu_acc_0_31017_37228);
  fu_acc_0_31017_37234 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_96_i0_fu_acc_0_31017_37234,
    in1 => out_const_36,
    in2 => out_extract_bit_expr_FU_65_i0_fu_acc_0_31017_37132,
    in3 => out_extract_bit_expr_FU_66_i0_fu_acc_0_31017_37135,
    in4 => out_extract_bit_expr_FU_67_i0_fu_acc_0_31017_37138,
    in5 => out_extract_bit_expr_FU_68_i0_fu_acc_0_31017_37141,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37237 : lut_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_97_i0_fu_acc_0_31017_37237,
    in1 => out_const_37,
    in2 => out_extract_bit_expr_FU_63_i0_fu_acc_0_31017_37126,
    in3 => out_extract_bit_expr_FU_64_i0_fu_acc_0_31017_37129,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919(0),
    in6 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in7 => out_lut_expr_FU_96_i0_fu_acc_0_31017_37234(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37240 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_98_i0_fu_acc_0_31017_37240,
    in1 => out_const_72,
    in2 => out_extract_bit_expr_FU_69_i0_fu_acc_0_31017_37144,
    in3 => out_extract_bit_expr_FU_70_i0_fu_acc_0_31017_37147,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in6 => out_lut_expr_FU_97_i0_fu_acc_0_31017_37237(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37243 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_99_i0_fu_acc_0_31017_37243,
    in1 => out_const_36,
    in2 => out_extract_bit_expr_FU_73_i0_fu_acc_0_31017_37156,
    in3 => out_extract_bit_expr_FU_74_i0_fu_acc_0_31017_37159,
    in4 => out_extract_bit_expr_FU_75_i0_fu_acc_0_31017_37162,
    in5 => out_extract_bit_expr_FU_76_i0_fu_acc_0_31017_37165,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37246 : lut_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_100_i0_fu_acc_0_31017_37246,
    in1 => out_const_37,
    in2 => out_extract_bit_expr_FU_71_i0_fu_acc_0_31017_37150,
    in3 => out_extract_bit_expr_FU_72_i0_fu_acc_0_31017_37153,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919(0),
    in6 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in7 => out_lut_expr_FU_99_i0_fu_acc_0_31017_37243(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37249 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_101_i0_fu_acc_0_31017_37249,
    in1 => out_const_72,
    in2 => out_extract_bit_expr_FU_77_i0_fu_acc_0_31017_37168,
    in3 => out_extract_bit_expr_FU_78_i0_fu_acc_0_31017_37171,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in6 => out_lut_expr_FU_100_i0_fu_acc_0_31017_37246(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37252 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_102_i0_fu_acc_0_31017_37252,
    in1 => out_const_36,
    in2 => out_extract_bit_expr_FU_81_i0_fu_acc_0_31017_37180,
    in3 => out_extract_bit_expr_FU_82_i0_fu_acc_0_31017_37183,
    in4 => out_extract_bit_expr_FU_83_i0_fu_acc_0_31017_37186,
    in5 => out_extract_bit_expr_FU_84_i0_fu_acc_0_31017_37189,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37255 : lut_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_103_i0_fu_acc_0_31017_37255,
    in1 => out_const_37,
    in2 => out_extract_bit_expr_FU_79_i0_fu_acc_0_31017_37174,
    in3 => out_extract_bit_expr_FU_80_i0_fu_acc_0_31017_37177,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919(0),
    in6 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in7 => out_lut_expr_FU_102_i0_fu_acc_0_31017_37252(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37258 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_104_i0_fu_acc_0_31017_37258,
    in1 => out_const_72,
    in2 => out_extract_bit_expr_FU_85_i0_fu_acc_0_31017_37192,
    in3 => out_extract_bit_expr_FU_86_i0_fu_acc_0_31017_37195,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in6 => out_lut_expr_FU_103_i0_fu_acc_0_31017_37255(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37261 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_105_i0_fu_acc_0_31017_37261,
    in1 => out_const_36,
    in2 => out_extract_bit_expr_FU_89_i0_fu_acc_0_31017_37204,
    in3 => out_extract_bit_expr_FU_90_i0_fu_acc_0_31017_37207,
    in4 => out_extract_bit_expr_FU_91_i0_fu_acc_0_31017_37210,
    in5 => out_extract_bit_expr_FU_92_i0_fu_acc_0_31017_37213,
    in6 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in7 => out_lut_expr_FU_24_i0_fu_acc_0_31017_36916(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37264 : lut_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_106_i0_fu_acc_0_31017_37264,
    in1 => out_const_37,
    in2 => out_extract_bit_expr_FU_87_i0_fu_acc_0_31017_37198,
    in3 => out_extract_bit_expr_FU_88_i0_fu_acc_0_31017_37201,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_25_i0_fu_acc_0_31017_36919(0),
    in6 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in7 => out_lut_expr_FU_105_i0_fu_acc_0_31017_37261(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37267 : lut_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_107_i0_fu_acc_0_31017_37267,
    in1 => out_const_72,
    in2 => out_extract_bit_expr_FU_93_i0_fu_acc_0_31017_37216,
    in3 => out_extract_bit_expr_FU_94_i0_fu_acc_0_31017_37219,
    in4 => out_lut_expr_FU_19_i0_fu_acc_0_31017_36835(0),
    in5 => out_lut_expr_FU_47_i0_fu_acc_0_31017_37009(0),
    in6 => out_lut_expr_FU_106_i0_fu_acc_0_31017_37264(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37270 : lut_expr_FU generic map(BITSIZE_in1=>59,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_108_i0_fu_acc_0_31017_37270,
    in1 => out_const_28,
    in2 => out_ui_eq_expr_FU_32_0_32_291_i4_fu_acc_0_31017_37123(0),
    in3 => out_lut_expr_FU_61_i0_fu_acc_0_31017_37054(0),
    in4 => out_lut_expr_FU_98_i0_fu_acc_0_31017_37240(0),
    in5 => out_lut_expr_FU_101_i0_fu_acc_0_31017_37249(0),
    in6 => out_lut_expr_FU_104_i0_fu_acc_0_31017_37258(0),
    in7 => out_lut_expr_FU_107_i0_fu_acc_0_31017_37267(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37273 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_109_i0_fu_acc_0_31017_37273,
    in1 => out_lut_expr_FU_108_i0_fu_acc_0_31017_37270);
  fu_acc_0_31017_37276 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>5,
    BITSIZE_out1=>5) port map (out1 => out_ui_bit_ior_expr_FU_0_8_8_285_i0_fu_acc_0_31017_37276,
    in1 => unsigned(out_UUdata_converter_FU_109_i0_fu_acc_0_31017_37273),
    in2 => out_ui_bit_ior_expr_FU_0_8_8_284_i0_fu_acc_0_31017_37231);
  fu_acc_0_31017_37279 : UIdata_converter_FU generic map(BITSIZE_in1=>5,
    BITSIZE_out1=>6) port map (out1 => out_UIdata_converter_FU_110_i0_fu_acc_0_31017_37279,
    in1 => out_ui_bit_ior_expr_FU_0_8_8_285_i0_fu_acc_0_31017_37276);
  fu_acc_0_31017_37282 : plus_expr_FU generic map(BITSIZE_in1=>6,
    BITSIZE_in2=>1,
    BITSIZE_out1=>7) port map (out1 => out_plus_expr_FU_8_0_8_261_i0_fu_acc_0_31017_37282,
    in1 => out_UIdata_converter_FU_110_i0_fu_acc_0_31017_37279,
    in2 => signed(out_const_15));
  fu_acc_0_31017_37285 : IIdata_converter_FU generic map(BITSIZE_in1=>7,
    BITSIZE_out1=>7) port map (out1 => out_IIdata_converter_FU_111_i0_fu_acc_0_31017_37285,
    in1 => out_plus_expr_FU_8_0_8_261_i0_fu_acc_0_31017_37282);
  fu_acc_0_31017_37288 : minus_expr_FU generic map(BITSIZE_in1=>9,
    BITSIZE_in2=>7,
    BITSIZE_out1=>9) port map (out1 => out_minus_expr_FU_0_8_8_257_i0_fu_acc_0_31017_37288,
    in1 => signed(out_const_7),
    in2 => out_IIdata_converter_FU_111_i0_fu_acc_0_31017_37285);
  fu_acc_0_31017_37291 : IUdata_converter_FU generic map(BITSIZE_in1=>9,
    BITSIZE_out1=>8) port map (out1 => out_IUdata_converter_FU_112_i0_fu_acc_0_31017_37291,
    in1 => out_minus_expr_FU_0_8_8_257_i0_fu_acc_0_31017_37288);
  fu_acc_0_31017_37294 : ui_lshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>6,
    BITSIZE_out1=>31,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_299_i0_fu_acc_0_31017_37294,
    in1 => out_IUdata_converter_FU_112_i0_fu_acc_0_31017_37291,
    in2 => out_const_9);
  fu_acc_0_31017_37297 : ui_rshift_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>5,
    BITSIZE_out1=>8,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_334_i0_fu_acc_0_31017_37297,
    in1 => out_ui_lshift_expr_FU_32_0_32_299_i0_fu_acc_0_31017_37294,
    in2 => out_const_40);
  fu_acc_0_31017_37300 : multi_read_cond_FU generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_multi_read_cond_FU_115_i0_fu_acc_0_31017_37300,
      in1(0 downto 0) => out_reg_12_reg_12);
  fu_acc_0_31017_37301 : ui_lshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>7,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in1 => unsigned(out_reg_14_reg_14),
    in2 => out_reg_15_reg_15);
  fu_acc_0_31017_37304 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3,
    BITSIZE_out1=>26,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_335_i0_fu_acc_0_31017_37304,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_43);
  fu_acc_0_31017_37307 : ui_plus_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>26,
    BITSIZE_out1=>26) port map (out1 => out_ui_plus_expr_FU_0_32_32_316_i0_fu_acc_0_31017_37307,
    in1 => unsigned(out_const_15),
    in2 => out_ui_rshift_expr_FU_32_0_32_335_i0_fu_acc_0_31017_37304);
  fu_acc_0_31017_37310 : ui_lshift_expr_FU generic map(BITSIZE_in1=>26,
    BITSIZE_in2=>3,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_300_i0_fu_acc_0_31017_37310,
    in1 => out_ui_plus_expr_FU_0_32_32_316_i0_fu_acc_0_31017_37307,
    in2 => out_const_43);
  fu_acc_0_31017_37313 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>4,
    BITSIZE_out1=>25,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_336_i0_fu_acc_0_31017_37313,
    in1 => out_ui_lshift_expr_FU_32_0_32_300_i0_fu_acc_0_31017_37310,
    in2 => out_const_13);
  fu_acc_0_31017_37316 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_240_i0_fu_acc_0_31017_37316,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_0);
  fu_acc_0_31017_37319 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_241_i0_fu_acc_0_31017_37319,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_15);
  fu_acc_0_31017_37322 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>2) port map (out1 => out_ui_extract_bit_expr_FU_242_i0_fu_acc_0_31017_37322,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_16);
  fu_acc_0_31017_37325 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>2) port map (out1 => out_ui_extract_bit_expr_FU_243_i0_fu_acc_0_31017_37325,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_42);
  fu_acc_0_31017_37328 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_ui_extract_bit_expr_FU_244_i0_fu_acc_0_31017_37328,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_17);
  fu_acc_0_31017_37331 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_ui_extract_bit_expr_FU_245_i0_fu_acc_0_31017_37331,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_33);
  fu_acc_0_31017_37334 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>3) port map (out1 => out_ui_extract_bit_expr_FU_246_i0_fu_acc_0_31017_37334,
    in1 => out_ui_lshift_expr_FU_32_32_32_303_i0_fu_acc_0_31017_37301,
    in2 => out_const_43);
  fu_acc_0_31017_37337 : lut_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_247_i0_fu_acc_0_31017_37337,
    in1 => out_const_25,
    in2 => out_ui_extract_bit_expr_FU_240_i0_fu_acc_0_31017_37316,
    in3 => out_ui_extract_bit_expr_FU_241_i0_fu_acc_0_31017_37319,
    in4 => out_ui_extract_bit_expr_FU_242_i0_fu_acc_0_31017_37322,
    in5 => out_ui_extract_bit_expr_FU_243_i0_fu_acc_0_31017_37325,
    in6 => out_ui_extract_bit_expr_FU_245_i0_fu_acc_0_31017_37331,
    in7 => out_ui_extract_bit_expr_FU_246_i0_fu_acc_0_31017_37334,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37340 : lut_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_248_i0_fu_acc_0_31017_37340,
    in1 => out_const_17,
    in2 => out_ui_extract_bit_expr_FU_244_i0_fu_acc_0_31017_37328,
    in3 => out_lut_expr_FU_247_i0_fu_acc_0_31017_37337(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37343 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_249_i0_fu_acc_0_31017_37343,
    in1 => unsigned(out_lut_expr_FU_248_i0_fu_acc_0_31017_37340));
  fu_acc_0_31017_37346 : bit_not_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>2) port map (out1 => out_bit_not_expr_FU_8_8_254_i0_fu_acc_0_31017_37346,
    in1 => out_UIdata_converter_FU_249_i0_fu_acc_0_31017_37343);
  fu_acc_0_31017_37349 : IUdata_converter_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>25) port map (out1 => out_IUdata_converter_FU_250_i0_fu_acc_0_31017_37349,
    in1 => out_bit_not_expr_FU_8_8_254_i0_fu_acc_0_31017_37346);
  fu_acc_0_31017_37352 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>25,
    BITSIZE_in2=>25,
    BITSIZE_out1=>25) port map (out1 => out_ui_bit_and_expr_FU_32_32_32_271_i0_fu_acc_0_31017_37352,
    in1 => out_ui_rshift_expr_FU_32_0_32_336_i0_fu_acc_0_31017_37313,
    in2 => out_IUdata_converter_FU_250_i0_fu_acc_0_31017_37349);
  fu_acc_0_31017_37355 : ui_eq_expr_FU generic map(BITSIZE_in1=>25,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_292_i0_fu_acc_0_31017_37355,
    in1 => out_ui_bit_and_expr_FU_32_32_32_271_i0_fu_acc_0_31017_37352,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37358 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>25,
    BITSIZE_in2=>31,
    BITSIZE_out1=>25) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_267_i0_fu_acc_0_31017_37358,
    in1 => out_ui_bit_and_expr_FU_32_32_32_271_i0_fu_acc_0_31017_37352,
    in2 => unsigned(out_const_75));
  fu_acc_0_31017_37361 : ui_bit_ior_concat_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>25,
    BITSIZE_in3=>5,
    BITSIZE_out1=>32,
    OFFSET_PARAMETER=>31) port map (out1 => out_ui_bit_ior_concat_expr_FU_276_i0_fu_acc_0_31017_37361,
    in1 => unsigned(out_reg_11_reg_11),
    in2 => out_ui_bit_and_expr_FU_32_0_32_267_i0_fu_acc_0_31017_37358,
    in3 => unsigned(out_const_62));
  fu_acc_0_31017_37364 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>9,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_334_i1_fu_acc_0_31017_37364,
    in1 => out_ui_bit_ior_concat_expr_FU_276_i0_fu_acc_0_31017_37361,
    in2 => out_const_40);
  fu_acc_0_31017_37367 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>23,
    BITSIZE_out1=>23) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_268_i0_fu_acc_0_31017_37367,
    in1 => out_ui_bit_ior_concat_expr_FU_276_i0_fu_acc_0_31017_37361,
    in2 => unsigned(out_const_73));
  fu_acc_0_31017_37370 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_in3=>8,
    BITSIZE_out1=>8) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i2_fu_acc_0_31017_37370,
    in1 => out_ui_eq_expr_FU_32_0_32_292_i0_fu_acc_0_31017_37355,
    in2 => unsigned(out_const_0),
    in3 => unsigned(out_reg_16_reg_16));
  fu_acc_0_31017_37373 : ui_lshift_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>5,
    BITSIZE_out1=>31,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_301_i0_fu_acc_0_31017_37373,
    in1 => out_ui_cond_expr_FU_8_8_8_8_289_i2_fu_acc_0_31017_37370,
    in2 => out_const_40);
  fu_acc_0_31017_37376 : ui_rshift_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>5,
    BITSIZE_out1=>8,
    PRECISION=>32) port map (out1 => out_ui_rshift_expr_FU_32_0_32_334_i2_fu_acc_0_31017_37376,
    in1 => out_ui_lshift_expr_FU_32_0_32_301_i0_fu_acc_0_31017_37373,
    in2 => out_const_40);
  fu_acc_0_31017_37379 : ui_plus_expr_FU generic map(BITSIZE_in1=>9,
    BITSIZE_in2=>8,
    BITSIZE_out1=>9) port map (out1 => out_ui_plus_expr_FU_8_8_8_319_i0_fu_acc_0_31017_37379,
    in1 => out_ui_rshift_expr_FU_32_0_32_334_i1_fu_acc_0_31017_37364,
    in2 => out_ui_rshift_expr_FU_32_0_32_334_i2_fu_acc_0_31017_37376);
  fu_acc_0_31017_37382 : ui_lshift_expr_FU generic map(BITSIZE_in1=>9,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    PRECISION=>32) port map (out1 => out_ui_lshift_expr_FU_32_0_32_301_i1_fu_acc_0_31017_37382,
    in1 => out_ui_plus_expr_FU_8_8_8_319_i0_fu_acc_0_31017_37379,
    in2 => out_const_40);
  fu_acc_0_31017_37385 : ui_bit_ior_concat_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>23,
    BITSIZE_in3=>5,
    BITSIZE_out1=>32,
    OFFSET_PARAMETER=>23) port map (out1 => out_ui_bit_ior_concat_expr_FU_277_i0_fu_acc_0_31017_37385,
    in1 => out_ui_lshift_expr_FU_32_0_32_301_i1_fu_acc_0_31017_37382,
    in2 => out_ui_bit_and_expr_FU_32_0_32_268_i0_fu_acc_0_31017_37367,
    in3 => unsigned(out_const_40));
  fu_acc_0_31017_37393 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>23,
    BITSIZE_out1=>23) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_269_i0_fu_acc_0_31017_37393,
    in1 => unsigned(out_UUdata_converter_FU_117_i0_fu_acc_0_31017_33178),
    in2 => unsigned(out_const_73));
  fu_acc_0_31017_37398 : ui_rshift_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>6,
    BITSIZE_out1=>8,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_337_i0_fu_acc_0_31017_37398,
    in1 => unsigned(out_UUdata_converter_FU_117_i0_fu_acc_0_31017_33178),
    in2 => out_const_9);
  fu_acc_0_31017_37401 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>8,
    BITSIZE_out1=>8) port map (out1 => out_ui_bit_and_expr_FU_8_0_8_275_i0_fu_acc_0_31017_37401,
    in1 => out_ui_rshift_expr_FU_32_0_32_337_i0_fu_acc_0_31017_37398,
    in2 => unsigned(out_const_65));
  fu_acc_0_31017_37404 : UUdata_converter_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>8) port map (out1 => out_UUdata_converter_FU_119_i0_fu_acc_0_31017_37404,
    in1 => std_logic_vector(out_ui_bit_and_expr_FU_8_0_8_275_i0_fu_acc_0_31017_37401));
  fu_acc_0_31017_37409 : ui_rshift_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>6,
    BITSIZE_out1=>8,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_337_i1_fu_acc_0_31017_37409,
    in1 => unsigned(out_UUdata_converter_FU_118_i0_fu_acc_0_31017_33181),
    in2 => out_const_9);
  fu_acc_0_31017_37414 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_in2=>8,
    BITSIZE_out1=>8) port map (out1 => out_ui_bit_and_expr_FU_0_8_8_265_i0_fu_acc_0_31017_37414,
    in1 => unsigned(out_const_65),
    in2 => out_ui_rshift_expr_FU_32_0_32_337_i1_fu_acc_0_31017_37409);
  fu_acc_0_31017_37417 : UUdata_converter_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>8) port map (out1 => out_UUdata_converter_FU_120_i0_fu_acc_0_31017_37417,
    in1 => std_logic_vector(out_ui_bit_and_expr_FU_0_8_8_265_i0_fu_acc_0_31017_37414));
  fu_acc_0_31017_37422 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>23,
    BITSIZE_out1=>23) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_269_i1_fu_acc_0_31017_37422,
    in1 => unsigned(out_UUdata_converter_FU_118_i0_fu_acc_0_31017_33181),
    in2 => unsigned(out_const_73));
  fu_acc_0_31017_37431 : lut_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_123_i0_fu_acc_0_31017_37431,
    in1 => out_const_43,
    in2 => out_reg_27_reg_27(0),
    in3 => out_ui_extract_bit_expr_FU_122_i0_fu_acc_0_31017_37955,
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37434 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_124_i0_fu_acc_0_31017_37434,
    in1 => out_lut_expr_FU_123_i0_fu_acc_0_31017_37431);
  fu_acc_0_31017_37437 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>6,
    BITSIZE_out1=>32,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_294_i1_fu_acc_0_31017_37437,
    in1 => unsigned(out_UUdata_converter_FU_124_i0_fu_acc_0_31017_37434),
    in2 => out_const_14);
  fu_acc_0_31017_37440 : ui_eq_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_293_i0_fu_acc_0_31017_37440,
    in1 => out_ui_bit_and_expr_FU_32_0_32_269_i0_fu_acc_0_31017_37393,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37473 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_135_i0_fu_acc_0_31017_37473,
    in1 => out_const_18,
    in2 => out_ui_eq_expr_FU_32_0_32_293_i0_fu_acc_0_31017_37440(0),
    in3 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37476 : ui_ne_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_ne_expr_FU_32_0_32_314_i0_fu_acc_0_31017_37476,
    in1 => out_ui_bit_and_expr_FU_32_0_32_269_i0_fu_acc_0_31017_37393,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37479 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_136_i0_fu_acc_0_31017_37479,
    in1 => out_const_18,
    in2 => out_ui_ne_expr_FU_32_0_32_314_i0_fu_acc_0_31017_37476(0),
    in3 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37482 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_in3=>1,
    BITSIZE_out1=>2) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i3_fu_acc_0_31017_37482,
    in1 => out_lut_expr_FU_136_i0_fu_acc_0_31017_37479,
    in2 => unsigned(out_const_42),
    in3 => unsigned(out_const_0));
  fu_acc_0_31017_37485 : ui_eq_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_293_i1_fu_acc_0_31017_37485,
    in1 => out_ui_bit_and_expr_FU_32_0_32_269_i1_fu_acc_0_31017_37422,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37518 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_147_i0_fu_acc_0_31017_37518,
    in1 => out_const_18,
    in2 => out_ui_eq_expr_FU_32_0_32_293_i1_fu_acc_0_31017_37485(0),
    in3 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37521 : ui_ne_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_ne_expr_FU_32_0_32_314_i1_fu_acc_0_31017_37521,
    in1 => out_ui_bit_and_expr_FU_32_0_32_269_i1_fu_acc_0_31017_37422,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37524 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_148_i0_fu_acc_0_31017_37524,
    in1 => out_const_18,
    in2 => out_ui_ne_expr_FU_32_0_32_314_i1_fu_acc_0_31017_37521(0),
    in3 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37527 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_in3=>1,
    BITSIZE_out1=>2) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i4_fu_acc_0_31017_37527,
    in1 => out_lut_expr_FU_148_i0_fu_acc_0_31017_37524,
    in2 => unsigned(out_const_42),
    in3 => unsigned(out_const_0));
  fu_acc_0_31017_37530 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>23,
    BITSIZE_out1=>24) port map (out1 => out_ui_bit_ior_expr_FU_0_32_32_278_i0_fu_acc_0_31017_37530,
    in1 => unsigned(out_const_23),
    in2 => out_ui_bit_and_expr_FU_32_0_32_269_i0_fu_acc_0_31017_37393);
  fu_acc_0_31017_37533 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>23,
    BITSIZE_out1=>24) port map (out1 => out_ui_bit_ior_expr_FU_0_32_32_278_i1_fu_acc_0_31017_37533,
    in1 => unsigned(out_const_23),
    in2 => out_ui_bit_and_expr_FU_32_0_32_269_i1_fu_acc_0_31017_37422);
  fu_acc_0_31017_37536 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>32,
    BITSIZE_out1=>24) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_270_i0_fu_acc_0_31017_37536,
    in1 => out_ui_bit_ior_expr_FU_0_32_32_278_i0_fu_acc_0_31017_37530,
    in2 => unsigned(out_const_76));
  fu_acc_0_31017_37539 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>32,
    BITSIZE_out1=>24) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_270_i1_fu_acc_0_31017_37539,
    in1 => out_ui_bit_ior_expr_FU_0_32_32_278_i1_fu_acc_0_31017_37533,
    in2 => unsigned(out_const_76));
  fu_acc_0_31017_37542 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_bit_ior_expr_FU_0_32_32_279_i0_fu_acc_0_31017_37542,
    in1 => unsigned(out_const_66),
    in2 => out_ui_lshift_expr_FU_32_0_32_294_i1_fu_acc_0_31017_37437);
  fu_acc_0_31017_37545 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_in3=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i5_fu_acc_0_31017_37545,
    in1 => out_lut_expr_FU_135_i0_fu_acc_0_31017_37473,
    in2 => unsigned(out_const_0),
    in3 => out_ui_cond_expr_FU_8_8_8_8_289_i3_fu_acc_0_31017_37482);
  fu_acc_0_31017_37548 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_149_i0_fu_acc_0_31017_37548,
    in1 => out_lut_expr_FU_135_i0_fu_acc_0_31017_37473);
  fu_acc_0_31017_37551 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_out1=>2,
    PRECISION=>8) port map (out1 => out_ui_lshift_expr_FU_8_0_8_312_i0_fu_acc_0_31017_37551,
    in1 => unsigned(out_UUdata_converter_FU_149_i0_fu_acc_0_31017_37548),
    in2 => out_const_15);
  fu_acc_0_31017_37581 : lut_expr_FU generic map(BITSIZE_in1=>12,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_159_i0_fu_acc_0_31017_37581,
    in1 => out_const_55,
    in2 => out_ui_extract_bit_expr_FU_154_i0_fu_acc_0_31017_38039,
    in3 => out_ui_extract_bit_expr_FU_155_i0_fu_acc_0_31017_38043,
    in4 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092(0),
    in5 => out_lut_expr_FU_158_i0_fu_acc_0_31017_38105(0),
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37584 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_160_i0_fu_acc_0_31017_37584,
    in1 => out_lut_expr_FU_159_i0_fu_acc_0_31017_37581);
  fu_acc_0_31017_37587 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_bit_ior_expr_FU_8_8_8_286_i0_fu_acc_0_31017_37587,
    in1 => out_ui_lshift_expr_FU_8_0_8_312_i0_fu_acc_0_31017_37551,
    in2 => out_ui_cond_expr_FU_8_8_8_8_289_i5_fu_acc_0_31017_37545);
  fu_acc_0_31017_37590 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_bit_ior_expr_FU_8_8_8_286_i1_fu_acc_0_31017_37590,
    in1 => unsigned(out_UUdata_converter_FU_160_i0_fu_acc_0_31017_37584),
    in2 => out_ui_bit_ior_expr_FU_8_8_8_286_i0_fu_acc_0_31017_37587);
  fu_acc_0_31017_37593 : ui_rshift_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>1,
    PRECISION=>8) port map (out1 => out_ui_rshift_expr_FU_8_0_8_344_i0_fu_acc_0_31017_37593,
    in1 => out_ui_bit_ior_expr_FU_8_8_8_286_i1_fu_acc_0_31017_37590,
    in2 => out_const_1);
  fu_acc_0_31017_37596 : UIdata_converter_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>3) port map (out1 => out_UIdata_converter_FU_161_i0_fu_acc_0_31017_37596,
    in1 => out_ui_bit_ior_expr_FU_8_8_8_286_i1_fu_acc_0_31017_37590);
  fu_acc_0_31017_37599 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_162_i0_fu_acc_0_31017_37599,
    in1 => out_ui_rshift_expr_FU_8_0_8_344_i0_fu_acc_0_31017_37593);
  fu_acc_0_31017_37602 : lut_expr_FU generic map(BITSIZE_in1=>61,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_163_i0_fu_acc_0_31017_37602,
    in1 => out_const_30,
    in2 => out_ui_eq_expr_FU_32_0_32_293_i0_fu_acc_0_31017_37440(0),
    in3 => out_ui_ne_expr_FU_32_0_32_314_i0_fu_acc_0_31017_37476(0),
    in4 => out_ui_extract_bit_expr_FU_154_i0_fu_acc_0_31017_38039,
    in5 => out_ui_extract_bit_expr_FU_155_i0_fu_acc_0_31017_38043,
    in6 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092(0),
    in7 => out_lut_expr_FU_158_i0_fu_acc_0_31017_38105(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37605 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_164_i0_fu_acc_0_31017_37605,
    in1 => out_lut_expr_FU_163_i0_fu_acc_0_31017_37602);
  fu_acc_0_31017_37608 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_165_i0_fu_acc_0_31017_37608,
    in1 => unsigned(out_UUdata_converter_FU_164_i0_fu_acc_0_31017_37605));
  fu_acc_0_31017_37611 : ui_ternary_plus_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>8,
    BITSIZE_in3=>8,
    BITSIZE_out1=>10) port map (out1 => out_ui_ternary_plus_expr_FU_0_16_16_16_345_i0_fu_acc_0_31017_37611,
    in1 => unsigned(out_const_74),
    in2 => unsigned(out_reg_20_reg_20),
    in3 => unsigned(out_UUdata_converter_FU_120_i0_fu_acc_0_31017_37417));
  fu_acc_0_31017_37614 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_in3=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_cond_expr_FU_8_8_8_8_289_i6_fu_acc_0_31017_37614,
    in1 => out_lut_expr_FU_147_i0_fu_acc_0_31017_37518,
    in2 => unsigned(out_const_0),
    in3 => out_ui_cond_expr_FU_8_8_8_8_289_i4_fu_acc_0_31017_37527);
  fu_acc_0_31017_37617 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_166_i0_fu_acc_0_31017_37617,
    in1 => out_lut_expr_FU_147_i0_fu_acc_0_31017_37518);
  fu_acc_0_31017_37620 : ui_lshift_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1,
    BITSIZE_out1=>2,
    PRECISION=>8) port map (out1 => out_ui_lshift_expr_FU_8_0_8_312_i1_fu_acc_0_31017_37620,
    in1 => unsigned(out_UUdata_converter_FU_166_i0_fu_acc_0_31017_37617),
    in2 => out_const_15);
  fu_acc_0_31017_37650 : lut_expr_FU generic map(BITSIZE_in1=>12,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_176_i0_fu_acc_0_31017_37650,
    in1 => out_const_55,
    in2 => out_ui_extract_bit_expr_FU_171_i0_fu_acc_0_31017_38071,
    in3 => out_ui_extract_bit_expr_FU_172_i0_fu_acc_0_31017_38075,
    in4 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100(0),
    in5 => out_lut_expr_FU_175_i0_fu_acc_0_31017_38110(0),
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37653 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_177_i0_fu_acc_0_31017_37653,
    in1 => out_lut_expr_FU_176_i0_fu_acc_0_31017_37650);
  fu_acc_0_31017_37656 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_bit_ior_expr_FU_8_8_8_286_i2_fu_acc_0_31017_37656,
    in1 => out_ui_lshift_expr_FU_8_0_8_312_i1_fu_acc_0_31017_37620,
    in2 => out_ui_cond_expr_FU_8_8_8_8_289_i6_fu_acc_0_31017_37614);
  fu_acc_0_31017_37659 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_ui_bit_ior_expr_FU_8_8_8_286_i3_fu_acc_0_31017_37659,
    in1 => unsigned(out_UUdata_converter_FU_177_i0_fu_acc_0_31017_37653),
    in2 => out_ui_bit_ior_expr_FU_8_8_8_286_i2_fu_acc_0_31017_37656);
  fu_acc_0_31017_37662 : ui_rshift_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>1,
    PRECISION=>8) port map (out1 => out_ui_rshift_expr_FU_8_0_8_344_i1_fu_acc_0_31017_37662,
    in1 => out_ui_bit_ior_expr_FU_8_8_8_286_i3_fu_acc_0_31017_37659,
    in2 => out_const_1);
  fu_acc_0_31017_37665 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>2,
    BITSIZE_out1=>1) port map (out1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in1 => out_ui_rshift_expr_FU_8_0_8_344_i1_fu_acc_0_31017_37662,
    in2 => out_ui_bit_ior_expr_FU_8_8_8_286_i3_fu_acc_0_31017_37659);
  fu_acc_0_31017_37668 : UIdata_converter_FU generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>3) port map (out1 => out_UIdata_converter_FU_178_i0_fu_acc_0_31017_37668,
    in1 => out_ui_bit_ior_expr_FU_8_8_8_286_i3_fu_acc_0_31017_37659);
  fu_acc_0_31017_37671 : bit_ior_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_in2=>2,
    BITSIZE_out1=>3) port map (out1 => out_bit_ior_expr_FU_8_8_8_253_i0_fu_acc_0_31017_37671,
    in1 => out_UIdata_converter_FU_178_i0_fu_acc_0_31017_37668,
    in2 => signed(out_reg_25_reg_25));
  fu_acc_0_31017_37674 : bit_and_expr_FU generic map(BITSIZE_in1=>3,
    BITSIZE_in2=>3,
    BITSIZE_out1=>2) port map (out1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in1 => out_bit_ior_expr_FU_8_8_8_253_i0_fu_acc_0_31017_37671,
    in2 => signed(out_reg_24_reg_24));
  fu_acc_0_31017_37677 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_179_i0_fu_acc_0_31017_37677,
    in1 => out_ui_rshift_expr_FU_8_0_8_344_i1_fu_acc_0_31017_37662);
  fu_acc_0_31017_37680 : bit_and_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in1 => signed(out_reg_26_reg_26),
    in2 => out_UIdata_converter_FU_179_i0_fu_acc_0_31017_37677);
  fu_acc_0_31017_37683 : lut_expr_FU generic map(BITSIZE_in1=>61,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_180_i0_fu_acc_0_31017_37683,
    in1 => out_const_30,
    in2 => out_ui_eq_expr_FU_32_0_32_293_i1_fu_acc_0_31017_37485(0),
    in3 => out_ui_ne_expr_FU_32_0_32_314_i1_fu_acc_0_31017_37521(0),
    in4 => out_ui_extract_bit_expr_FU_171_i0_fu_acc_0_31017_38071,
    in5 => out_ui_extract_bit_expr_FU_172_i0_fu_acc_0_31017_38075,
    in6 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100(0),
    in7 => out_lut_expr_FU_175_i0_fu_acc_0_31017_38110(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37686 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_181_i0_fu_acc_0_31017_37686,
    in1 => out_lut_expr_FU_180_i0_fu_acc_0_31017_37683);
  fu_acc_0_31017_37689 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_182_i0_fu_acc_0_31017_37689,
    in1 => unsigned(out_UUdata_converter_FU_181_i0_fu_acc_0_31017_37686));
  fu_acc_0_31017_37692 : bit_and_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>2,
    BITSIZE_out1=>2) port map (out1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in1 => out_UIdata_converter_FU_182_i0_fu_acc_0_31017_37689,
    in2 => signed(out_reg_25_reg_25));
  fu_acc_0_31017_37695 : ui_mult_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>24,
    BITSIZE_out1=>48,
    PIPE_PARAMETER=>0) port map (out1 => out_ui_mult_expr_FU_32_32_32_0_313_i0_fu_acc_0_31017_37695,
    clock => clock,
    in1 => unsigned(out_reg_23_reg_23),
    in2 => out_ui_bit_and_expr_FU_32_0_32_270_i1_fu_acc_0_31017_37539);
  fu_acc_0_31017_37698 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_in2=>6) port map (out1 => out_ui_extract_bit_expr_FU_183_i0_fu_acc_0_31017_37698,
    in1 => out_ui_mult_expr_FU_32_32_32_0_313_i0_fu_acc_0_31017_37695,
    in2 => out_const_41);
  fu_acc_0_31017_37701 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_184_i0_fu_acc_0_31017_37701,
    in1(0) => out_ui_extract_bit_expr_FU_183_i0_fu_acc_0_31017_37698);
  fu_acc_0_31017_37704 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_185_i0_fu_acc_0_31017_37704,
    in1 => out_UUdata_converter_FU_184_i0_fu_acc_0_31017_37701);
  fu_acc_0_31017_37707 : ui_plus_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>10,
    BITSIZE_out1=>10) port map (out1 => out_ui_plus_expr_FU_16_16_16_317_i0_fu_acc_0_31017_37707,
    in1 => unsigned(out_reg_34_reg_34),
    in2 => unsigned(out_reg_32_reg_32));
  fu_acc_0_31017_37710 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_in2=>6) port map (out1 => out_ui_extract_bit_expr_FU_186_i0_fu_acc_0_31017_37710,
    in1 => out_ui_mult_expr_FU_32_32_32_0_313_i0_fu_acc_0_31017_37695,
    in2 => out_const_41);
  fu_acc_0_31017_37713 : lut_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_187_i0_fu_acc_0_31017_37713,
    in1 => out_const_15,
    in2 => out_ui_extract_bit_expr_FU_186_i0_fu_acc_0_31017_37710,
    in3 => '0',
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37716 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_188_i0_fu_acc_0_31017_37716,
    in1 => out_lut_expr_FU_187_i0_fu_acc_0_31017_37713);
  fu_acc_0_31017_37719 : UIdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>2) port map (out1 => out_UIdata_converter_FU_189_i0_fu_acc_0_31017_37719,
    in1 => unsigned(out_UUdata_converter_FU_188_i0_fu_acc_0_31017_37716));
  fu_acc_0_31017_37722 : ui_lshift_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_in2=>2,
    BITSIZE_out1=>47,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_64_64_64_306_i0_fu_acc_0_31017_37722,
    in1 => unsigned(out_reg_33_reg_33),
    in2 => out_reg_35_reg_35);
  fu_acc_0_31017_37725 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>47,
    BITSIZE_in2=>47,
    BITSIZE_out1=>47) port map (out1 => out_ui_bit_and_expr_FU_0_64_64_263_i0_fu_acc_0_31017_37725,
    in1 => unsigned(out_const_78),
    in2 => out_ui_lshift_expr_FU_64_64_64_306_i0_fu_acc_0_31017_37722);
  fu_acc_0_31017_37728 : ui_lshift_expr_FU generic map(BITSIZE_in1=>47,
    BITSIZE_in2=>2,
    BITSIZE_out1=>48,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_64_0_64_304_i0_fu_acc_0_31017_37728,
    in1 => out_ui_bit_and_expr_FU_0_64_64_263_i0_fu_acc_0_31017_37725,
    in2 => out_const_1);
  fu_acc_0_31017_37731 : UUdata_converter_FU generic map(BITSIZE_in1=>10,
    BITSIZE_out1=>10) port map (out1 => out_UUdata_converter_FU_190_i0_fu_acc_0_31017_37731,
    in1 => std_logic_vector(out_ui_plus_expr_FU_16_16_16_317_i0_fu_acc_0_31017_37707));
  fu_acc_0_31017_37734 : ui_lshift_expr_FU generic map(BITSIZE_in1=>10,
    BITSIZE_in2=>6,
    BITSIZE_out1=>33,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_64_0_64_305_i0_fu_acc_0_31017_37734,
    in1 => unsigned(out_UUdata_converter_FU_190_i0_fu_acc_0_31017_37731),
    in2 => out_const_9);
  fu_acc_0_31017_37737 : ui_rshift_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_in2=>6,
    BITSIZE_out1=>23,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_64_0_64_340_i0_fu_acc_0_31017_37737,
    in1 => out_ui_lshift_expr_FU_64_0_64_304_i0_fu_acc_0_31017_37728,
    in2 => out_const_12);
  fu_acc_0_31017_37740 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>23,
    BITSIZE_out1=>23) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_269_i2_fu_acc_0_31017_37740,
    in1 => out_ui_rshift_expr_FU_64_0_64_340_i0_fu_acc_0_31017_37737,
    in2 => unsigned(out_const_73));
  fu_acc_0_31017_37743 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>23,
    BITSIZE_out1=>33) port map (out1 => out_ui_bit_ior_expr_FU_0_64_64_281_i0_fu_acc_0_31017_37743,
    in1 => out_ui_lshift_expr_FU_64_0_64_305_i0_fu_acc_0_31017_37734,
    in2 => out_ui_bit_and_expr_FU_32_0_32_269_i2_fu_acc_0_31017_37740);
  fu_acc_0_31017_37746 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>33,
    BITSIZE_out1=>33) port map (out1 => out_ui_bit_and_expr_FU_0_64_64_264_i0_fu_acc_0_31017_37746,
    in1 => unsigned(out_const_77),
    in2 => out_ui_bit_ior_expr_FU_0_64_64_281_i0_fu_acc_0_31017_37743);
  fu_acc_0_31017_37749 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>10,
    BITSIZE_in2=>4) port map (out1 => out_ui_extract_bit_expr_FU_191_i0_fu_acc_0_31017_37749,
    in1 => out_ui_plus_expr_FU_16_16_16_317_i0_fu_acc_0_31017_37707,
    in2 => out_const_31);
  fu_acc_0_31017_37752 : ui_rshift_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_in2=>1,
    BITSIZE_out1=>23,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_64_0_64_341_i0_fu_acc_0_31017_37752,
    in1 => out_ui_lshift_expr_FU_64_0_64_304_i0_fu_acc_0_31017_37728,
    in2 => out_const_15);
  fu_acc_0_31017_37755 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>23,
    BITSIZE_out1=>23) port map (out1 => out_ui_bit_and_expr_FU_32_0_32_269_i3_fu_acc_0_31017_37755,
    in1 => out_ui_rshift_expr_FU_64_0_64_341_i0_fu_acc_0_31017_37752,
    in2 => unsigned(out_const_73));
  fu_acc_0_31017_37758 : ui_lshift_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>24,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_298_i2_fu_acc_0_31017_37758,
    in1 => out_ui_bit_and_expr_FU_32_0_32_269_i3_fu_acc_0_31017_37755,
    in2 => out_const_15);
  fu_acc_0_31017_37761 : ui_rshift_expr_FU generic map(BITSIZE_in1=>24,
    BITSIZE_in2=>1,
    BITSIZE_out1=>23,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_332_i3_fu_acc_0_31017_37761,
    in1 => out_ui_lshift_expr_FU_32_0_32_298_i2_fu_acc_0_31017_37758,
    in2 => out_const_15);
  fu_acc_0_31017_37764 : ui_ne_expr_FU generic map(BITSIZE_in1=>23,
    BITSIZE_in2=>1,
    BITSIZE_out1=>1) port map (out1 => out_ui_ne_expr_FU_32_0_32_315_i0_fu_acc_0_31017_37764,
    in1 => out_ui_rshift_expr_FU_32_0_32_332_i3_fu_acc_0_31017_37761,
    in2 => unsigned(out_const_0));
  fu_acc_0_31017_37767 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>47,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_192_i0_fu_acc_0_31017_37767,
    in1 => out_ui_lshift_expr_FU_64_64_64_306_i0_fu_acc_0_31017_37722,
    in2 => out_const_44);
  fu_acc_0_31017_37770 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>47,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_193_i0_fu_acc_0_31017_37770,
    in1 => out_ui_lshift_expr_FU_64_64_64_306_i0_fu_acc_0_31017_37722,
    in2 => out_const_40);
  fu_acc_0_31017_37773 : lut_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_194_i0_fu_acc_0_31017_37773,
    in1 => out_const_53,
    in2 => out_ui_ne_expr_FU_32_0_32_315_i0_fu_acc_0_31017_37764(0),
    in3 => out_ui_extract_bit_expr_FU_192_i0_fu_acc_0_31017_37767,
    in4 => out_ui_extract_bit_expr_FU_193_i0_fu_acc_0_31017_37770,
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37776 : UUdata_converter_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_UUdata_converter_FU_195_i0_fu_acc_0_31017_37776,
    in1 => out_lut_expr_FU_194_i0_fu_acc_0_31017_37773);
  fu_acc_0_31017_37779 : ui_plus_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>1,
    BITSIZE_out1=>33) port map (out1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in1 => out_ui_bit_and_expr_FU_0_64_64_264_i0_fu_acc_0_31017_37746,
    in2 => unsigned(out_UUdata_converter_FU_195_i0_fu_acc_0_31017_37776));
  fu_acc_0_31017_37782 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>10,
    BITSIZE_in2=>4) port map (out1 => out_ui_extract_bit_expr_FU_196_i0_fu_acc_0_31017_37782,
    in1 => out_ui_plus_expr_FU_16_16_16_317_i0_fu_acc_0_31017_37707,
    in2 => out_const_31);
  fu_acc_0_31017_37785 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>6) port map (out1 => out_ui_extract_bit_expr_FU_197_i0_fu_acc_0_31017_37785,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_20);
  fu_acc_0_31017_37788 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_198_i0_fu_acc_0_31017_37788,
    in1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in2 => out_const_0);
  fu_acc_0_31017_37791 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_199_i0_fu_acc_0_31017_37791,
    in1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in2 => out_const_0);
  fu_acc_0_31017_37794 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_200_i0_fu_acc_0_31017_37794,
    in1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in2 => out_const_0);
  fu_acc_0_31017_37797 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_201_i0_fu_acc_0_31017_37797,
    in1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in2 => out_const_0);
  fu_acc_0_31017_37803 : lut_expr_FU generic map(BITSIZE_in1=>17,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_203_i0_fu_acc_0_31017_37803,
    in1 => out_const_22,
    in2 => out_extract_bit_expr_FU_198_i0_fu_acc_0_31017_37788,
    in3 => out_extract_bit_expr_FU_199_i0_fu_acc_0_31017_37791,
    in4 => out_ui_extract_bit_expr_FU_200_i0_fu_acc_0_31017_37794,
    in5 => out_extract_bit_expr_FU_201_i0_fu_acc_0_31017_37797,
    in6 => out_lut_expr_FU_202_i0_fu_acc_0_31017_38117(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37806 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_204_i0_fu_acc_0_31017_37806,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_40);
  fu_acc_0_31017_37809 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_205_i0_fu_acc_0_31017_37809,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_44);
  fu_acc_0_31017_37812 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_206_i0_fu_acc_0_31017_37812,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_45);
  fu_acc_0_31017_37815 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_207_i0_fu_acc_0_31017_37815,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_48);
  fu_acc_0_31017_37818 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_208_i0_fu_acc_0_31017_37818,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_49);
  fu_acc_0_31017_37821 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_209_i0_fu_acc_0_31017_37821,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_52);
  fu_acc_0_31017_37824 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_210_i0_fu_acc_0_31017_37824,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_57);
  fu_acc_0_31017_37827 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_211_i0_fu_acc_0_31017_37827,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_60);
  fu_acc_0_31017_37830 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>33,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_212_i0_fu_acc_0_31017_37830,
    in1 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779,
    in2 => out_const_62);
  fu_acc_0_31017_37833 : ui_bit_and_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>33,
    BITSIZE_out1=>31) port map (out1 => out_ui_bit_and_expr_FU_0_32_32_262_i0_fu_acc_0_31017_37833,
    in1 => unsigned(out_const_75),
    in2 => out_ui_plus_expr_FU_32_32_32_318_i0_fu_acc_0_31017_37779);
  fu_acc_0_31017_37836 : ui_bit_ior_expr_FU generic map(BITSIZE_in1=>31,
    BITSIZE_in2=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_bit_ior_expr_FU_0_32_32_280_i0_fu_acc_0_31017_37836,
    in1 => out_ui_bit_and_expr_FU_0_32_32_262_i0_fu_acc_0_31017_37833,
    in2 => unsigned(out_reg_30_reg_30));
  fu_acc_0_31017_37839 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_213_i0_fu_acc_0_31017_37839,
    in1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in2 => out_const_0);
  fu_acc_0_31017_37842 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_214_i0_fu_acc_0_31017_37842,
    in1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in2 => out_const_0);
  fu_acc_0_31017_37845 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_215_i0_fu_acc_0_31017_37845,
    in1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in2 => out_const_0);
  fu_acc_0_31017_37848 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_216_i0_fu_acc_0_31017_37848,
    in1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in2 => out_const_0);
  fu_acc_0_31017_37851 : lut_expr_FU generic map(BITSIZE_in1=>17,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_217_i0_fu_acc_0_31017_37851,
    in1 => out_const_71,
    in2 => out_extract_bit_expr_FU_213_i0_fu_acc_0_31017_37839,
    in3 => out_extract_bit_expr_FU_214_i0_fu_acc_0_31017_37842,
    in4 => out_ui_extract_bit_expr_FU_215_i0_fu_acc_0_31017_37845,
    in5 => out_extract_bit_expr_FU_216_i0_fu_acc_0_31017_37848,
    in6 => out_lut_expr_FU_202_i0_fu_acc_0_31017_38117(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37854 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_218_i0_fu_acc_0_31017_37854,
    in1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in2 => out_const_0);
  fu_acc_0_31017_37857 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_219_i0_fu_acc_0_31017_37857,
    in1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in2 => out_const_0);
  fu_acc_0_31017_37860 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_220_i0_fu_acc_0_31017_37860,
    in1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in2 => out_const_0);
  fu_acc_0_31017_37863 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_221_i0_fu_acc_0_31017_37863,
    in1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in2 => out_const_0);
  fu_acc_0_31017_37878 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_226_i0_fu_acc_0_31017_37878,
    in1 => out_const_18,
    in2 => out_reg_46_reg_46(0),
    in3 => out_lut_expr_FU_225_i0_fu_acc_0_31017_38132(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37881 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_227_i0_fu_acc_0_31017_37881,
    in1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in2 => out_const_0);
  fu_acc_0_31017_37884 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_228_i0_fu_acc_0_31017_37884,
    in1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in2 => out_const_0);
  fu_acc_0_31017_37887 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_229_i0_fu_acc_0_31017_37887,
    in1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in2 => out_const_0);
  fu_acc_0_31017_37890 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_230_i0_fu_acc_0_31017_37890,
    in1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in2 => out_const_0);
  fu_acc_0_31017_37896 : lut_expr_FU generic map(BITSIZE_in1=>4,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_232_i0_fu_acc_0_31017_37896,
    in1 => out_const_18,
    in2 => out_reg_46_reg_46(0),
    in3 => out_lut_expr_FU_231_i0_fu_acc_0_31017_38137(0),
    in4 => '0',
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37899 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>32,
    BITSIZE_in3=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i4_fu_acc_0_31017_37899,
    in1 => out_lut_expr_FU_232_i0_fu_acc_0_31017_37896,
    in2 => out_ui_bit_ior_expr_FU_0_32_32_280_i0_fu_acc_0_31017_37836,
    in3 => unsigned(out_reg_30_reg_30));
  fu_acc_0_31017_37902 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>32,
    BITSIZE_in3=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i5_fu_acc_0_31017_37902,
    in1 => out_lut_expr_FU_226_i0_fu_acc_0_31017_37878,
    in2 => unsigned(out_reg_31_reg_31),
    in3 => out_ui_cond_expr_FU_32_32_32_32_288_i4_fu_acc_0_31017_37899);
  fu_acc_0_31017_37905 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>10,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_338_i0_fu_acc_0_31017_37905,
    in1 => out_ui_lshift_expr_FU_32_0_32_294_i1_fu_acc_0_31017_37437,
    in2 => out_const_39);
  fu_acc_0_31017_37908 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>10,
    BITSIZE_in3=>10,
    BITSIZE_out1=>10) port map (out1 => out_ui_cond_expr_FU_16_16_16_16_287_i0_fu_acc_0_31017_37908,
    in1 => out_lut_expr_FU_203_i0_fu_acc_0_31017_37803,
    in2 => out_ui_rshift_expr_FU_32_0_32_338_i0_fu_acc_0_31017_37905,
    in3 => unsigned(out_const_67));
  fu_acc_0_31017_37911 : ui_lshift_expr_FU generic map(BITSIZE_in1=>10,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_302_i0_fu_acc_0_31017_37911,
    in1 => out_ui_cond_expr_FU_16_16_16_16_287_i0_fu_acc_0_31017_37908,
    in2 => out_const_39);
  fu_acc_0_31017_37914 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_233_i0_fu_acc_0_31017_37914,
    in1 => out_bit_and_expr_FU_8_8_8_252_i1_fu_acc_0_31017_37680,
    in2 => out_const_0);
  fu_acc_0_31017_37917 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_234_i0_fu_acc_0_31017_37917,
    in1 => out_bit_and_expr_FU_8_8_8_252_i2_fu_acc_0_31017_37692,
    in2 => out_const_0);
  fu_acc_0_31017_37920 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>1) port map (out1 => out_ui_extract_bit_expr_FU_235_i0_fu_acc_0_31017_37920,
    in1 => out_ui_bit_and_expr_FU_1_1_1_266_i0_fu_acc_0_31017_37665,
    in2 => out_const_0);
  fu_acc_0_31017_37923 : extract_bit_expr_FU generic map(BITSIZE_in1=>2,
    BITSIZE_in2=>1) port map (out1 => out_extract_bit_expr_FU_236_i0_fu_acc_0_31017_37923,
    in1 => out_bit_and_expr_FU_8_8_8_252_i0_fu_acc_0_31017_37674,
    in2 => out_const_0);
  fu_acc_0_31017_37926 : lut_expr_FU generic map(BITSIZE_in1=>17,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_237_i0_fu_acc_0_31017_37926,
    in1 => out_const_70,
    in2 => out_extract_bit_expr_FU_233_i0_fu_acc_0_31017_37914,
    in3 => out_extract_bit_expr_FU_234_i0_fu_acc_0_31017_37917,
    in4 => out_ui_extract_bit_expr_FU_235_i0_fu_acc_0_31017_37920,
    in5 => out_extract_bit_expr_FU_236_i0_fu_acc_0_31017_37923,
    in6 => out_lut_expr_FU_202_i0_fu_acc_0_31017_38117(0),
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_37929 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>10,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_339_i0_fu_acc_0_31017_37929,
    in1 => out_ui_lshift_expr_FU_32_0_32_302_i0_fu_acc_0_31017_37911,
    in2 => out_const_39);
  fu_acc_0_31017_37932 : ui_rshift_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5,
    BITSIZE_out1=>10,
    PRECISION=>64) port map (out1 => out_ui_rshift_expr_FU_32_0_32_338_i1_fu_acc_0_31017_37932,
    in1 => out_ui_bit_ior_expr_FU_0_32_32_279_i0_fu_acc_0_31017_37542,
    in2 => out_const_39);
  fu_acc_0_31017_37935 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>10,
    BITSIZE_in3=>10,
    BITSIZE_out1=>10) port map (out1 => out_ui_cond_expr_FU_16_16_16_16_287_i1_fu_acc_0_31017_37935,
    in1 => out_lut_expr_FU_237_i0_fu_acc_0_31017_37926,
    in2 => out_ui_rshift_expr_FU_32_0_32_339_i0_fu_acc_0_31017_37929,
    in3 => out_ui_rshift_expr_FU_32_0_32_338_i1_fu_acc_0_31017_37932);
  fu_acc_0_31017_37938 : ui_lshift_expr_FU generic map(BITSIZE_in1=>10,
    BITSIZE_in2=>5,
    BITSIZE_out1=>32,
    PRECISION=>64) port map (out1 => out_ui_lshift_expr_FU_32_0_32_302_i1_fu_acc_0_31017_37938,
    in1 => out_ui_cond_expr_FU_16_16_16_16_287_i1_fu_acc_0_31017_37935,
    in2 => out_const_39);
  fu_acc_0_31017_37941 : ui_cond_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_in2=>32,
    BITSIZE_in3=>32,
    BITSIZE_out1=>32) port map (out1 => out_ui_cond_expr_FU_32_32_32_32_288_i6_fu_acc_0_31017_37941,
    in1 => out_reg_36_reg_36,
    in2 => unsigned(out_reg_45_reg_45),
    in3 => out_ui_cond_expr_FU_32_32_32_32_288_i5_fu_acc_0_31017_37902);
  fu_acc_0_31017_37951 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_121_i0_fu_acc_0_31017_37951,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_62);
  fu_acc_0_31017_37955 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_122_i0_fu_acc_0_31017_37955,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_62);
  fu_acc_0_31017_37959 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_125_i0_fu_acc_0_31017_37959,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_40);
  fu_acc_0_31017_37963 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_126_i0_fu_acc_0_31017_37963,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_44);
  fu_acc_0_31017_37967 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_127_i0_fu_acc_0_31017_37967,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_45);
  fu_acc_0_31017_37971 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_128_i0_fu_acc_0_31017_37971,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_48);
  fu_acc_0_31017_37975 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_129_i0_fu_acc_0_31017_37975,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_49);
  fu_acc_0_31017_37979 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_130_i0_fu_acc_0_31017_37979,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_52);
  fu_acc_0_31017_37983 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_131_i0_fu_acc_0_31017_37983,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_57);
  fu_acc_0_31017_37987 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_132_i0_fu_acc_0_31017_37987,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_60);
  fu_acc_0_31017_37991 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_137_i0_fu_acc_0_31017_37991,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_40);
  fu_acc_0_31017_37995 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_138_i0_fu_acc_0_31017_37995,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_44);
  fu_acc_0_31017_37999 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_139_i0_fu_acc_0_31017_37999,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_45);
  fu_acc_0_31017_38003 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_140_i0_fu_acc_0_31017_38003,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_48);
  fu_acc_0_31017_38007 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_141_i0_fu_acc_0_31017_38007,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_49);
  fu_acc_0_31017_38011 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_142_i0_fu_acc_0_31017_38011,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_52);
  fu_acc_0_31017_38015 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_143_i0_fu_acc_0_31017_38015,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_57);
  fu_acc_0_31017_38019 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_144_i0_fu_acc_0_31017_38019,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_60);
  fu_acc_0_31017_38023 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_150_i0_fu_acc_0_31017_38023,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_49);
  fu_acc_0_31017_38027 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_151_i0_fu_acc_0_31017_38027,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_52);
  fu_acc_0_31017_38031 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_152_i0_fu_acc_0_31017_38031,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_57);
  fu_acc_0_31017_38035 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_153_i0_fu_acc_0_31017_38035,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_60);
  fu_acc_0_31017_38039 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_154_i0_fu_acc_0_31017_38039,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_40);
  fu_acc_0_31017_38043 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_155_i0_fu_acc_0_31017_38043,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_44);
  fu_acc_0_31017_38047 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_156_i0_fu_acc_0_31017_38047,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_45);
  fu_acc_0_31017_38051 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_157_i0_fu_acc_0_31017_38051,
    in1 => unsigned(out_reg_13_reg_13),
    in2 => out_const_48);
  fu_acc_0_31017_38055 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_167_i0_fu_acc_0_31017_38055,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_49);
  fu_acc_0_31017_38059 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_168_i0_fu_acc_0_31017_38059,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_52);
  fu_acc_0_31017_38063 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_169_i0_fu_acc_0_31017_38063,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_57);
  fu_acc_0_31017_38067 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_170_i0_fu_acc_0_31017_38067,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_60);
  fu_acc_0_31017_38071 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_171_i0_fu_acc_0_31017_38071,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_40);
  fu_acc_0_31017_38075 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_172_i0_fu_acc_0_31017_38075,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_44);
  fu_acc_0_31017_38079 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_173_i0_fu_acc_0_31017_38079,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_45);
  fu_acc_0_31017_38083 : ui_extract_bit_expr_FU generic map(BITSIZE_in1=>32,
    BITSIZE_in2=>5) port map (out1 => out_ui_extract_bit_expr_FU_174_i0_fu_acc_0_31017_38083,
    in1 => unsigned(out_reg_29_reg_29),
    in2 => out_const_48);
  fu_acc_0_31017_38089 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_133_i0_fu_acc_0_31017_38089,
    in1 => out_const_26,
    in2 => out_ui_extract_bit_expr_FU_125_i0_fu_acc_0_31017_37959,
    in3 => out_ui_extract_bit_expr_FU_126_i0_fu_acc_0_31017_37963,
    in4 => out_ui_extract_bit_expr_FU_127_i0_fu_acc_0_31017_37967,
    in5 => out_ui_extract_bit_expr_FU_128_i0_fu_acc_0_31017_37971,
    in6 => out_ui_extract_bit_expr_FU_131_i0_fu_acc_0_31017_37983,
    in7 => out_ui_extract_bit_expr_FU_132_i0_fu_acc_0_31017_37987,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38092 : lut_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092,
    in1 => out_const_21,
    in2 => out_ui_extract_bit_expr_FU_129_i0_fu_acc_0_31017_37975,
    in3 => out_ui_extract_bit_expr_FU_130_i0_fu_acc_0_31017_37979,
    in4 => out_lut_expr_FU_133_i0_fu_acc_0_31017_38089(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38097 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_145_i0_fu_acc_0_31017_38097,
    in1 => out_const_26,
    in2 => out_ui_extract_bit_expr_FU_137_i0_fu_acc_0_31017_37991,
    in3 => out_ui_extract_bit_expr_FU_138_i0_fu_acc_0_31017_37995,
    in4 => out_ui_extract_bit_expr_FU_139_i0_fu_acc_0_31017_37999,
    in5 => out_ui_extract_bit_expr_FU_140_i0_fu_acc_0_31017_38003,
    in6 => out_ui_extract_bit_expr_FU_143_i0_fu_acc_0_31017_38015,
    in7 => out_ui_extract_bit_expr_FU_144_i0_fu_acc_0_31017_38019,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38100 : lut_expr_FU generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100,
    in1 => out_const_21,
    in2 => out_ui_extract_bit_expr_FU_141_i0_fu_acc_0_31017_38007,
    in3 => out_ui_extract_bit_expr_FU_142_i0_fu_acc_0_31017_38011,
    in4 => out_lut_expr_FU_145_i0_fu_acc_0_31017_38097(0),
    in5 => '0',
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38105 : lut_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_158_i0_fu_acc_0_31017_38105,
    in1 => out_const_15,
    in2 => out_ui_extract_bit_expr_FU_150_i0_fu_acc_0_31017_38023,
    in3 => out_ui_extract_bit_expr_FU_151_i0_fu_acc_0_31017_38027,
    in4 => out_ui_extract_bit_expr_FU_152_i0_fu_acc_0_31017_38031,
    in5 => out_ui_extract_bit_expr_FU_153_i0_fu_acc_0_31017_38035,
    in6 => out_ui_extract_bit_expr_FU_156_i0_fu_acc_0_31017_38047,
    in7 => out_ui_extract_bit_expr_FU_157_i0_fu_acc_0_31017_38051,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38110 : lut_expr_FU generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_175_i0_fu_acc_0_31017_38110,
    in1 => out_const_15,
    in2 => out_ui_extract_bit_expr_FU_167_i0_fu_acc_0_31017_38055,
    in3 => out_ui_extract_bit_expr_FU_168_i0_fu_acc_0_31017_38059,
    in4 => out_ui_extract_bit_expr_FU_169_i0_fu_acc_0_31017_38063,
    in5 => out_ui_extract_bit_expr_FU_170_i0_fu_acc_0_31017_38067,
    in6 => out_ui_extract_bit_expr_FU_173_i0_fu_acc_0_31017_38079,
    in7 => out_ui_extract_bit_expr_FU_174_i0_fu_acc_0_31017_38083,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38117 : lut_expr_FU generic map(BITSIZE_in1=>49,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_202_i0_fu_acc_0_31017_38117,
    in1 => out_const_27,
    in2 => out_reg_21_reg_21(0),
    in3 => out_reg_22_reg_22(0),
    in4 => out_ui_eq_expr_FU_32_0_32_293_i1_fu_acc_0_31017_37485(0),
    in5 => out_ui_ne_expr_FU_32_0_32_314_i1_fu_acc_0_31017_37521(0),
    in6 => out_reg_28_reg_28(0),
    in7 => out_lut_expr_FU_146_i0_fu_acc_0_31017_38100(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38122 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_222_i0_fu_acc_0_31017_38122,
    in1 => out_const_26,
    in2 => out_ui_extract_bit_expr_FU_204_i0_fu_acc_0_31017_37806,
    in3 => out_ui_extract_bit_expr_FU_205_i0_fu_acc_0_31017_37809,
    in4 => out_ui_extract_bit_expr_FU_206_i0_fu_acc_0_31017_37812,
    in5 => out_ui_extract_bit_expr_FU_207_i0_fu_acc_0_31017_37815,
    in6 => out_ui_extract_bit_expr_FU_210_i0_fu_acc_0_31017_37824,
    in7 => out_ui_extract_bit_expr_FU_211_i0_fu_acc_0_31017_37827,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38125 : lut_expr_FU generic map(BITSIZE_in1=>11,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_223_i0_fu_acc_0_31017_38125,
    in1 => out_const_56,
    in2 => out_ui_extract_bit_expr_FU_208_i0_fu_acc_0_31017_37818,
    in3 => out_ui_extract_bit_expr_FU_209_i0_fu_acc_0_31017_37821,
    in4 => out_ui_extract_bit_expr_FU_212_i0_fu_acc_0_31017_37830,
    in5 => out_lut_expr_FU_222_i0_fu_acc_0_31017_38122(0),
    in6 => '0',
    in7 => '0',
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38128 : lut_expr_FU generic map(BITSIZE_in1=>56,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_224_i0_fu_acc_0_31017_38128,
    in1 => out_const_54,
    in2 => out_ui_ne_expr_FU_32_0_32_315_i0_fu_acc_0_31017_37764(0),
    in3 => out_ui_extract_bit_expr_FU_192_i0_fu_acc_0_31017_37767,
    in4 => out_ui_extract_bit_expr_FU_193_i0_fu_acc_0_31017_37770,
    in5 => out_ui_extract_bit_expr_FU_196_i0_fu_acc_0_31017_37782,
    in6 => out_ui_extract_bit_expr_FU_197_i0_fu_acc_0_31017_37785,
    in7 => out_ui_extract_bit_expr_FU_191_i0_fu_acc_0_31017_37749,
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38132 : lut_expr_FU generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_225_i0_fu_acc_0_31017_38132,
    in1 => out_const_68,
    in2 => out_reg_37_reg_37(0),
    in3 => out_reg_38_reg_38(0),
    in4 => out_reg_39_reg_39(0),
    in5 => out_reg_40_reg_40(0),
    in6 => out_lut_expr_FU_223_i0_fu_acc_0_31017_38125(0),
    in7 => out_lut_expr_FU_224_i0_fu_acc_0_31017_38128(0),
    in8 => '0',
    in9 => '0');
  fu_acc_0_31017_38137 : lut_expr_FU generic map(BITSIZE_in1=>64,
    BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_231_i0_fu_acc_0_31017_38137,
    in1 => out_const_69,
    in2 => out_reg_41_reg_41(0),
    in3 => out_reg_42_reg_42(0),
    in4 => out_reg_43_reg_43(0),
    in5 => out_reg_44_reg_44(0),
    in6 => out_lut_expr_FU_223_i0_fu_acc_0_31017_38125(0),
    in7 => out_lut_expr_FU_224_i0_fu_acc_0_31017_38128(0),
    in8 => '0',
    in9 => '0');
  s_MEMORY_CTRL_D21_251_i00 <= selector_IN_UNBOUNDED_acc_0_31017_31056 or selector_IN_UNBOUNDED_acc_0_31017_31057 or selector_IN_UNBOUNDED_acc_0_31017_31059 or selector_IN_UNBOUNDED_acc_0_31017_31060 or selector_IN_UNBOUNDED_acc_0_31017_31061 or selector_IN_UNBOUNDED_acc_0_31017_31063 or selector_IN_UNBOUNDED_acc_0_31017_31065 or selector_IN_UNBOUNDED_acc_0_31017_31066 or selector_IN_UNBOUNDED_acc_0_31017_31068;
  reg_0 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_0_reg_0,
    clock => clock,
    reset => reset,
    in1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    wenable => wrenable_reg_0);
  reg_1 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_1_reg_1,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_3_i0_fu_acc_0_31017_31446,
    wenable => wrenable_reg_1);
  reg_10 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_10_reg_10,
    clock => clock,
    reset => reset,
    in1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    wenable => wrenable_reg_10);
  reg_11 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_11_reg_11,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_lshift_expr_FU_32_0_32_295_i0_fu_acc_0_31017_36829),
    wenable => wrenable_reg_11);
  reg_12 : register_SE generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_12_reg_12,
    clock => clock,
    reset => reset,
    in1 => out_lut_expr_FU_20_i0_fu_acc_0_31017_36838,
    wenable => wrenable_reg_12);
  reg_13 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_13_reg_13,
    clock => clock,
    reset => reset,
    in1 => out_MUX_550_reg_13_0_0_0,
    wenable => wrenable_reg_13);
  reg_14 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_14_reg_14,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_cond_expr_FU_32_32_32_32_288_i0_fu_acc_0_31017_36847),
    wenable => wrenable_reg_14);
  reg_15 : register_SE generic map(BITSIZE_in1=>7,
    BITSIZE_out1=>7) port map (out1 => out_reg_15_reg_15,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_IIdata_converter_FU_111_i0_fu_acc_0_31017_37285),
    wenable => wrenable_reg_15);
  reg_16 : register_SE generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>8) port map (out1 => out_reg_16_reg_16,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_rshift_expr_FU_32_0_32_334_i0_fu_acc_0_31017_37297),
    wenable => wrenable_reg_16);
  reg_17 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_17_reg_17,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_mult_expr_FU_32_32_32_0_258_i0_fu_acc_0_31017_31062),
    wenable => wrenable_reg_17);
  reg_18 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_18_reg_18,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_plus_expr_FU_32_32_32_260_i0_fu_acc_0_31017_31058),
    wenable => wrenable_reg_18);
  reg_19 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_19_reg_19,
    clock => clock,
    reset => reset,
    in1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    wenable => wrenable_reg_19);
  reg_2 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_2_reg_2,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_5_i0_fu_acc_0_31017_31466,
    wenable => wrenable_reg_2);
  reg_20 : register_SE generic map(BITSIZE_in1=>8,
    BITSIZE_out1=>8) port map (out1 => out_reg_20_reg_20,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_119_i0_fu_acc_0_31017_37404,
    wenable => wrenable_reg_20);
  reg_21 : register_SE generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_21_reg_21,
    clock => clock,
    reset => reset,
    in1 => out_ui_eq_expr_FU_32_0_32_293_i0_fu_acc_0_31017_37440,
    wenable => wrenable_reg_21);
  reg_22 : register_SE generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_22_reg_22,
    clock => clock,
    reset => reset,
    in1 => out_ui_ne_expr_FU_32_0_32_314_i0_fu_acc_0_31017_37476,
    wenable => wrenable_reg_22);
  reg_23 : register_SE generic map(BITSIZE_in1=>24,
    BITSIZE_out1=>24) port map (out1 => out_reg_23_reg_23,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_bit_and_expr_FU_32_0_32_270_i0_fu_acc_0_31017_37536),
    wenable => wrenable_reg_23);
  reg_24 : register_SE generic map(BITSIZE_in1=>3,
    BITSIZE_out1=>3) port map (out1 => out_reg_24_reg_24,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_UIdata_converter_FU_161_i0_fu_acc_0_31017_37596),
    wenable => wrenable_reg_24);
  reg_25 : register_SE generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>2) port map (out1 => out_reg_25_reg_25,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_UIdata_converter_FU_162_i0_fu_acc_0_31017_37599),
    wenable => wrenable_reg_25);
  reg_26 : register_SE generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>2) port map (out1 => out_reg_26_reg_26,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_UIdata_converter_FU_165_i0_fu_acc_0_31017_37608),
    wenable => wrenable_reg_26);
  reg_27 : register_SE generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_27_reg_27,
    clock => clock,
    reset => reset,
    in1(0) => out_ui_extract_bit_expr_FU_121_i0_fu_acc_0_31017_37951,
    wenable => wrenable_reg_27);
  reg_28 : register_SE generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_28_reg_28,
    clock => clock,
    reset => reset,
    in1 => out_lut_expr_FU_134_i0_fu_acc_0_31017_38092,
    wenable => wrenable_reg_28);
  reg_29 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_29_reg_29,
    clock => clock,
    reset => reset,
    in1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    wenable => wrenable_reg_29);
  reg_3 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_3_reg_3,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_7_i0_fu_acc_0_31017_31479,
    wenable => wrenable_reg_3);
  reg_30 : register_STD generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_30_reg_30,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_lshift_expr_FU_32_0_32_294_i1_fu_acc_0_31017_37437),
    wenable => wrenable_reg_30);
  reg_31 : register_STD generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_31_reg_31,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_bit_ior_expr_FU_0_32_32_279_i0_fu_acc_0_31017_37542),
    wenable => wrenable_reg_31);
  reg_32 : register_STD generic map(BITSIZE_in1=>10,
    BITSIZE_out1=>10) port map (out1 => out_reg_32_reg_32,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_ternary_plus_expr_FU_0_16_16_16_345_i0_fu_acc_0_31017_37611),
    wenable => wrenable_reg_32);
  reg_33 : register_STD generic map(BITSIZE_in1=>48,
    BITSIZE_out1=>48) port map (out1 => out_reg_33_reg_33,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_mult_expr_FU_32_32_32_0_313_i0_fu_acc_0_31017_37695),
    wenable => wrenable_reg_33);
  reg_34 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_34_reg_34,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_185_i0_fu_acc_0_31017_37704,
    wenable => wrenable_reg_34);
  reg_35 : register_STD generic map(BITSIZE_in1=>2,
    BITSIZE_out1=>2) port map (out1 => out_reg_35_reg_35,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_UIdata_converter_FU_189_i0_fu_acc_0_31017_37719),
    wenable => wrenable_reg_35);
  reg_36 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_36_reg_36,
    clock => clock,
    reset => reset,
    in1 => out_lut_expr_FU_217_i0_fu_acc_0_31017_37851,
    wenable => wrenable_reg_36);
  reg_37 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_37_reg_37,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_218_i0_fu_acc_0_31017_37854,
    wenable => wrenable_reg_37);
  reg_38 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_38_reg_38,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_219_i0_fu_acc_0_31017_37857,
    wenable => wrenable_reg_38);
  reg_39 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_39_reg_39,
    clock => clock,
    reset => reset,
    in1(0) => out_ui_extract_bit_expr_FU_220_i0_fu_acc_0_31017_37860,
    wenable => wrenable_reg_39);
  reg_4 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_4_reg_4,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_320_i0_fu_acc_0_31017_31501),
    wenable => wrenable_reg_4);
  reg_40 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_40_reg_40,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_221_i0_fu_acc_0_31017_37863,
    wenable => wrenable_reg_40);
  reg_41 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_41_reg_41,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_227_i0_fu_acc_0_31017_37881,
    wenable => wrenable_reg_41);
  reg_42 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_42_reg_42,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_228_i0_fu_acc_0_31017_37884,
    wenable => wrenable_reg_42);
  reg_43 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_43_reg_43,
    clock => clock,
    reset => reset,
    in1(0) => out_ui_extract_bit_expr_FU_229_i0_fu_acc_0_31017_37887,
    wenable => wrenable_reg_43);
  reg_44 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_44_reg_44,
    clock => clock,
    reset => reset,
    in1(0) => out_extract_bit_expr_FU_230_i0_fu_acc_0_31017_37890,
    wenable => wrenable_reg_44);
  reg_45 : register_STD generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_45_reg_45,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_lshift_expr_FU_32_0_32_302_i1_fu_acc_0_31017_37938),
    wenable => wrenable_reg_45);
  reg_46 : register_STD generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => out_reg_46_reg_46,
    clock => clock,
    reset => reset,
    in1 => out_lut_expr_FU_202_i0_fu_acc_0_31017_38117,
    wenable => wrenable_reg_46);
  reg_47 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_47_reg_47,
    clock => clock,
    reset => reset,
    in1 => out_UUdata_converter_FU_238_i0_fu_acc_0_31017_33175,
    wenable => wrenable_reg_47);
  reg_5 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_5_reg_5,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_320_i1_fu_acc_0_31017_31514),
    wenable => wrenable_reg_5);
  reg_6 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_6_reg_6,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_320_i2_fu_acc_0_31017_31527),
    wenable => wrenable_reg_6);
  reg_7 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_7_reg_7,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_322_i0_fu_acc_0_31017_31625),
    wenable => wrenable_reg_7);
  reg_8 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_8_reg_8,
    clock => clock,
    reset => reset,
    in1 => std_logic_vector(out_ui_pointer_plus_expr_FU_32_0_32_321_i2_fu_acc_0_31017_31632),
    wenable => wrenable_reg_8);
  reg_9 : register_SE generic map(BITSIZE_in1=>32,
    BITSIZE_out1=>32) port map (out1 => out_reg_9_reg_9,
    clock => clock,
    reset => reset,
    in1 => out_MEMORY_CTRL_D21_251_i0_MEMORY_CTRL_D21_251_i0,
    wenable => wrenable_reg_9);
  -- io-signal post fix
  Mout_oe_ram <= \sig_out_bus_mergerMout_oe_ram3_\(0);
  Mout_we_ram <= \sig_out_bus_mergerMout_we_ram4_\(0);
  Mout_addr_ram <= \sig_out_bus_mergerMout_addr_ram1_\;
  Mout_Wdata_ram <= \sig_out_bus_mergerMout_Wdata_ram0_\;
  Mout_data_ram_size <= \sig_out_bus_mergerMout_data_ram_size2_\;
  OUT_MULTIIF_acc_0_31017_37300 <= out_multi_read_cond_FU_115_i0_fu_acc_0_31017_37300;
  OUT_UNBOUNDED_acc_0_31017_31056 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31057 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31059 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31060 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31061 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31063 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31065 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31066 <= s_done_MEMORY_CTRL_D21_251_i0;
  OUT_UNBOUNDED_acc_0_31017_31068 <= s_done_MEMORY_CTRL_D21_251_i0;

end datapath_acc_0_arch;

-- FSM based controller description for acc_0
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity controller_acc_0 is 
port (
  -- IN
  OUT_MULTIIF_acc_0_31017_37300 : in std_logic_vector(0 downto 0);
  OUT_UNBOUNDED_acc_0_31017_31056 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31057 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31059 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31060 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31061 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31063 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31065 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31066 : in std_logic;
  OUT_UNBOUNDED_acc_0_31017_31068 : in std_logic;
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  -- OUT
  done_port : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31056 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31057 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31059 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31060 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31061 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31063 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31065 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31066 : out std_logic;
  selector_IN_UNBOUNDED_acc_0_31017_31068 : out std_logic;
  fuselector_MEMORY_CTRL_D21_251_i0_LOAD : out std_logic;
  fuselector_MEMORY_CTRL_D21_251_i0_STORE : out std_logic;
  selector_MUX_550_reg_13_0_0_0 : out std_logic;
  selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : out std_logic;
  selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : out std_logic;
  selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : out std_logic;
  wrenable_reg_0 : out std_logic;
  wrenable_reg_1 : out std_logic;
  wrenable_reg_10 : out std_logic;
  wrenable_reg_11 : out std_logic;
  wrenable_reg_12 : out std_logic;
  wrenable_reg_13 : out std_logic;
  wrenable_reg_14 : out std_logic;
  wrenable_reg_15 : out std_logic;
  wrenable_reg_16 : out std_logic;
  wrenable_reg_17 : out std_logic;
  wrenable_reg_18 : out std_logic;
  wrenable_reg_19 : out std_logic;
  wrenable_reg_2 : out std_logic;
  wrenable_reg_20 : out std_logic;
  wrenable_reg_21 : out std_logic;
  wrenable_reg_22 : out std_logic;
  wrenable_reg_23 : out std_logic;
  wrenable_reg_24 : out std_logic;
  wrenable_reg_25 : out std_logic;
  wrenable_reg_26 : out std_logic;
  wrenable_reg_27 : out std_logic;
  wrenable_reg_28 : out std_logic;
  wrenable_reg_29 : out std_logic;
  wrenable_reg_3 : out std_logic;
  wrenable_reg_30 : out std_logic;
  wrenable_reg_31 : out std_logic;
  wrenable_reg_32 : out std_logic;
  wrenable_reg_33 : out std_logic;
  wrenable_reg_34 : out std_logic;
  wrenable_reg_35 : out std_logic;
  wrenable_reg_36 : out std_logic;
  wrenable_reg_37 : out std_logic;
  wrenable_reg_38 : out std_logic;
  wrenable_reg_39 : out std_logic;
  wrenable_reg_4 : out std_logic;
  wrenable_reg_40 : out std_logic;
  wrenable_reg_41 : out std_logic;
  wrenable_reg_42 : out std_logic;
  wrenable_reg_43 : out std_logic;
  wrenable_reg_44 : out std_logic;
  wrenable_reg_45 : out std_logic;
  wrenable_reg_46 : out std_logic;
  wrenable_reg_47 : out std_logic;
  wrenable_reg_5 : out std_logic;
  wrenable_reg_6 : out std_logic;
  wrenable_reg_7 : out std_logic;
  wrenable_reg_8 : out std_logic;
  wrenable_reg_9 : out std_logic

);
end controller_acc_0;

architecture controller_acc_0_arch of controller_acc_0 is
  -- define the states of FSM model
  constant S_0: std_logic_vector(22 downto 0) := "00000000000000000000001";
  constant S_1: std_logic_vector(22 downto 0) := "00000000000000000000010";
  constant S_2: std_logic_vector(22 downto 0) := "00000000000000000000100";
  constant S_3: std_logic_vector(22 downto 0) := "00000000000000000001000";
  constant S_4: std_logic_vector(22 downto 0) := "00000000000000000010000";
  constant S_5: std_logic_vector(22 downto 0) := "00000000000000000100000";
  constant S_6: std_logic_vector(22 downto 0) := "00000000000000001000000";
  constant S_7: std_logic_vector(22 downto 0) := "00000000000000010000000";
  constant S_8: std_logic_vector(22 downto 0) := "00000000000000100000000";
  constant S_9: std_logic_vector(22 downto 0) := "00000000000001000000000";
  constant S_10: std_logic_vector(22 downto 0) := "00000000000010000000000";
  constant S_11: std_logic_vector(22 downto 0) := "00000000000100000000000";
  constant S_12: std_logic_vector(22 downto 0) := "00000000001000000000000";
  constant S_22: std_logic_vector(22 downto 0) := "10000000000000000000000";
  constant S_13: std_logic_vector(22 downto 0) := "00000000010000000000000";
  constant S_14: std_logic_vector(22 downto 0) := "00000000100000000000000";
  constant S_15: std_logic_vector(22 downto 0) := "00000001000000000000000";
  constant S_16: std_logic_vector(22 downto 0) := "00000010000000000000000";
  constant S_17: std_logic_vector(22 downto 0) := "00000100000000000000000";
  constant S_18: std_logic_vector(22 downto 0) := "00001000000000000000000";
  constant S_19: std_logic_vector(22 downto 0) := "00010000000000000000000";
  constant S_20: std_logic_vector(22 downto 0) := "00100000000000000000000";
  constant S_21: std_logic_vector(22 downto 0) := "01000000000000000000000";
  signal present_state : std_logic_vector(22 downto 0) := S_0;
  signal next_state : std_logic_vector(22 downto 0);
begin
  -- concurrent process#1: state registers
  state_reg: process(clock)
  begin
    if (clock'event and clock='1') then
      if (reset='0') then
        present_state <= S_0;
      else
        present_state <= next_state;
      end if;
    end if;
  end process;
  -- concurrent process#0: combinational logic
  comb_logic0: process(present_state, OUT_MULTIIF_acc_0_31017_37300, OUT_UNBOUNDED_acc_0_31017_31056, OUT_UNBOUNDED_acc_0_31017_31057, OUT_UNBOUNDED_acc_0_31017_31059, OUT_UNBOUNDED_acc_0_31017_31060, OUT_UNBOUNDED_acc_0_31017_31061, OUT_UNBOUNDED_acc_0_31017_31063, OUT_UNBOUNDED_acc_0_31017_31065, OUT_UNBOUNDED_acc_0_31017_31066, OUT_UNBOUNDED_acc_0_31017_31068, start_port)
  begin
    done_port <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31056 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31057 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31059 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31060 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31061 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31063 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31065 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31066 <= '0';
    selector_IN_UNBOUNDED_acc_0_31017_31068 <= '0';
    fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '0';
    fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '0';
    selector_MUX_550_reg_13_0_0_0 <= '0';
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 <= '0';
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 <= '0';
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '0';
    wrenable_reg_0 <= '0';
    wrenable_reg_1 <= '0';
    wrenable_reg_10 <= '0';
    wrenable_reg_11 <= '0';
    wrenable_reg_12 <= '0';
    wrenable_reg_13 <= '0';
    wrenable_reg_14 <= '0';
    wrenable_reg_15 <= '0';
    wrenable_reg_16 <= '0';
    wrenable_reg_17 <= '0';
    wrenable_reg_18 <= '0';
    wrenable_reg_19 <= '0';
    wrenable_reg_2 <= '0';
    wrenable_reg_20 <= '0';
    wrenable_reg_21 <= '0';
    wrenable_reg_22 <= '0';
    wrenable_reg_23 <= '0';
    wrenable_reg_24 <= '0';
    wrenable_reg_25 <= '0';
    wrenable_reg_26 <= '0';
    wrenable_reg_27 <= '0';
    wrenable_reg_28 <= '0';
    wrenable_reg_29 <= '0';
    wrenable_reg_3 <= '0';
    wrenable_reg_30 <= '0';
    wrenable_reg_31 <= '0';
    wrenable_reg_32 <= '0';
    wrenable_reg_33 <= '0';
    wrenable_reg_34 <= '0';
    wrenable_reg_35 <= '0';
    wrenable_reg_36 <= '0';
    wrenable_reg_37 <= '0';
    wrenable_reg_38 <= '0';
    wrenable_reg_39 <= '0';
    wrenable_reg_4 <= '0';
    wrenable_reg_40 <= '0';
    wrenable_reg_41 <= '0';
    wrenable_reg_42 <= '0';
    wrenable_reg_43 <= '0';
    wrenable_reg_44 <= '0';
    wrenable_reg_45 <= '0';
    wrenable_reg_46 <= '0';
    wrenable_reg_47 <= '0';
    wrenable_reg_5 <= '0';
    wrenable_reg_6 <= '0';
    wrenable_reg_7 <= '0';
    wrenable_reg_8 <= '0';
    wrenable_reg_9 <= '0';
    next_state <= S_0;
    case present_state is
      when S_0 =>
        if(start_port /= '1') then
          selector_MUX_550_reg_13_0_0_0 <= 'X';
          selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 <= 'X';
          selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 <= 'X';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= 'X';
          wrenable_reg_0 <= 'X';
          wrenable_reg_1 <= 'X';
          wrenable_reg_10 <= 'X';
          wrenable_reg_11 <= 'X';
          wrenable_reg_12 <= 'X';
          wrenable_reg_13 <= 'X';
          wrenable_reg_14 <= 'X';
          wrenable_reg_15 <= 'X';
          wrenable_reg_16 <= 'X';
          wrenable_reg_17 <= 'X';
          wrenable_reg_18 <= 'X';
          wrenable_reg_19 <= 'X';
          wrenable_reg_2 <= 'X';
          wrenable_reg_20 <= 'X';
          wrenable_reg_21 <= 'X';
          wrenable_reg_22 <= 'X';
          wrenable_reg_23 <= 'X';
          wrenable_reg_24 <= 'X';
          wrenable_reg_25 <= 'X';
          wrenable_reg_26 <= 'X';
          wrenable_reg_27 <= 'X';
          wrenable_reg_28 <= 'X';
          wrenable_reg_29 <= 'X';
          wrenable_reg_3 <= 'X';
          wrenable_reg_30 <= 'X';
          wrenable_reg_31 <= 'X';
          wrenable_reg_32 <= 'X';
          wrenable_reg_33 <= 'X';
          wrenable_reg_34 <= 'X';
          wrenable_reg_35 <= 'X';
          wrenable_reg_36 <= 'X';
          wrenable_reg_37 <= 'X';
          wrenable_reg_38 <= 'X';
          wrenable_reg_39 <= 'X';
          wrenable_reg_4 <= 'X';
          wrenable_reg_40 <= 'X';
          wrenable_reg_41 <= 'X';
          wrenable_reg_42 <= 'X';
          wrenable_reg_43 <= 'X';
          wrenable_reg_44 <= 'X';
          wrenable_reg_45 <= 'X';
          wrenable_reg_46 <= 'X';
          wrenable_reg_47 <= 'X';
          wrenable_reg_5 <= 'X';
          wrenable_reg_6 <= 'X';
          wrenable_reg_7 <= 'X';
          wrenable_reg_8 <= 'X';
          wrenable_reg_9 <= 'X';
          next_state <= S_0;
        else
          selector_IN_UNBOUNDED_acc_0_31017_31056 <= '1';
          fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
          selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 <= '1';
          wrenable_reg_0 <= OUT_UNBOUNDED_acc_0_31017_31056;
          wrenable_reg_1 <= '1';
          wrenable_reg_2 <= '1';
          wrenable_reg_3 <= '1';
          wrenable_reg_4 <= '1';
          wrenable_reg_5 <= '1';
          wrenable_reg_6 <= '1';
          wrenable_reg_7 <= '1';
          wrenable_reg_8 <= '1';
          if (OUT_UNBOUNDED_acc_0_31017_31056 = '0') then
            next_state <= S_1;
          else
            next_state <= S_2;
          end if;
        end if;
      when S_1 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 <= '1';
        wrenable_reg_0 <= OUT_UNBOUNDED_acc_0_31017_31056;
        if (OUT_UNBOUNDED_acc_0_31017_31056 = '0') then
          next_state <= S_1;
        else
          next_state <= S_2;
        end if;
      when S_2 =>
        selector_IN_UNBOUNDED_acc_0_31017_31060 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_9 <= OUT_UNBOUNDED_acc_0_31017_31060;
        if (OUT_UNBOUNDED_acc_0_31017_31060 = '0') then
          next_state <= S_3;
        else
          next_state <= S_4;
        end if;
      when S_3 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_9 <= OUT_UNBOUNDED_acc_0_31017_31060;
        if (OUT_UNBOUNDED_acc_0_31017_31060 = '0') then
          next_state <= S_3;
        else
          next_state <= S_4;
        end if;
      when S_4 =>
        selector_IN_UNBOUNDED_acc_0_31017_31061 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        wrenable_reg_10 <= OUT_UNBOUNDED_acc_0_31017_31061;
        wrenable_reg_11 <= '1';
        wrenable_reg_12 <= '1';
        wrenable_reg_13 <= '1';
        wrenable_reg_14 <= '1';
        wrenable_reg_15 <= '1';
        wrenable_reg_16 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31061 = '0') then
          next_state <= S_5;
        else
          next_state <= S_6;
        end if;
      when S_5 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        wrenable_reg_10 <= OUT_UNBOUNDED_acc_0_31017_31061;
        if (OUT_UNBOUNDED_acc_0_31017_31061 = '0') then
          next_state <= S_5;
        else
          next_state <= S_6;
        end if;
      when S_6 =>
        selector_IN_UNBOUNDED_acc_0_31017_31057 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_17 <= '1';
        wrenable_reg_9 <= OUT_UNBOUNDED_acc_0_31017_31057;
        if (OUT_UNBOUNDED_acc_0_31017_31057 = '0') then
          next_state <= S_7;
        else
          next_state <= S_8;
        end if;
      when S_7 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_9 <= OUT_UNBOUNDED_acc_0_31017_31057;
        if (OUT_UNBOUNDED_acc_0_31017_31057 = '0') then
          next_state <= S_7;
        else
          next_state <= S_8;
        end if;
      when S_8 =>
        selector_IN_UNBOUNDED_acc_0_31017_31063 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 <= '1';
        wrenable_reg_18 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31063 = '0') then
          next_state <= S_9;
        else
          next_state <= S_10;
        end if;
      when S_9 =>
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31063 = '0') then
          next_state <= S_9;
        else
          next_state <= S_10;
        end if;
      when S_10 =>
        selector_IN_UNBOUNDED_acc_0_31017_31059 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31059 = '0') then
          next_state <= S_11;
        else
          next_state <= S_12;
        end if;
      when S_11 =>
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31059 = '0') then
          next_state <= S_11;
        else
          next_state <= S_12;
        end if;
      when S_12 =>
        if (OUT_MULTIIF_acc_0_31017_37300(0) = '1') then
          next_state <= S_22;
        else
          next_state <= S_13;
        end if;
      when S_22 =>
        selector_MUX_550_reg_13_0_0_0 <= '1';
        wrenable_reg_13 <= '1';
        next_state <= S_13;
      when S_13 =>
        selector_IN_UNBOUNDED_acc_0_31017_31065 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= '1';
        wrenable_reg_19 <= OUT_UNBOUNDED_acc_0_31017_31065;
        wrenable_reg_20 <= '1';
        wrenable_reg_21 <= '1';
        wrenable_reg_22 <= '1';
        wrenable_reg_23 <= '1';
        wrenable_reg_24 <= '1';
        wrenable_reg_25 <= '1';
        wrenable_reg_26 <= '1';
        wrenable_reg_27 <= '1';
        wrenable_reg_28 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31065 = '0') then
          next_state <= S_14;
        else
          next_state <= S_15;
        end if;
      when S_14 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= '1';
        wrenable_reg_19 <= OUT_UNBOUNDED_acc_0_31017_31065;
        if (OUT_UNBOUNDED_acc_0_31017_31065 = '0') then
          next_state <= S_14;
        else
          next_state <= S_15;
        end if;
      when S_15 =>
        selector_IN_UNBOUNDED_acc_0_31017_31066 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_29 <= OUT_UNBOUNDED_acc_0_31017_31066;
        if (OUT_UNBOUNDED_acc_0_31017_31066 = '0') then
          next_state <= S_16;
        else
          next_state <= S_17;
        end if;
      when S_16 =>
        fuselector_MEMORY_CTRL_D21_251_i0_LOAD <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= '1';
        wrenable_reg_29 <= OUT_UNBOUNDED_acc_0_31017_31066;
        if (OUT_UNBOUNDED_acc_0_31017_31066 = '0') then
          next_state <= S_16;
        else
          next_state <= S_17;
        end if;
      when S_17 =>
        wrenable_reg_30 <= '1';
        wrenable_reg_31 <= '1';
        wrenable_reg_32 <= '1';
        wrenable_reg_33 <= '1';
        wrenable_reg_34 <= '1';
        wrenable_reg_35 <= '1';
        wrenable_reg_36 <= '1';
        wrenable_reg_37 <= '1';
        wrenable_reg_38 <= '1';
        wrenable_reg_39 <= '1';
        wrenable_reg_40 <= '1';
        wrenable_reg_41 <= '1';
        wrenable_reg_42 <= '1';
        wrenable_reg_43 <= '1';
        wrenable_reg_44 <= '1';
        wrenable_reg_45 <= '1';
        wrenable_reg_46 <= '1';
        next_state <= S_18;
      when S_18 =>
        wrenable_reg_47 <= '1';
        next_state <= S_19;
      when S_19 =>
        selector_IN_UNBOUNDED_acc_0_31017_31068 <= '1';
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31068 = '0') then
          next_state <= S_20;
        else
          next_state <= S_21;
          done_port <= '1';
        end if;
      when S_20 =>
        fuselector_MEMORY_CTRL_D21_251_i0_STORE <= '1';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 <= '1';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= '1';
        if (OUT_UNBOUNDED_acc_0_31017_31068 = '0') then
          next_state <= S_20;
        else
          next_state <= S_21;
          done_port <= '1';
        end if;
      when S_21 =>
        next_state <= S_0;
      when others =>
        selector_MUX_550_reg_13_0_0_0 <= 'X';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 <= 'X';
        selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 <= 'X';
        selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 <= 'X';
        wrenable_reg_0 <= 'X';
        wrenable_reg_1 <= 'X';
        wrenable_reg_10 <= 'X';
        wrenable_reg_11 <= 'X';
        wrenable_reg_12 <= 'X';
        wrenable_reg_13 <= 'X';
        wrenable_reg_14 <= 'X';
        wrenable_reg_15 <= 'X';
        wrenable_reg_16 <= 'X';
        wrenable_reg_17 <= 'X';
        wrenable_reg_18 <= 'X';
        wrenable_reg_19 <= 'X';
        wrenable_reg_2 <= 'X';
        wrenable_reg_20 <= 'X';
        wrenable_reg_21 <= 'X';
        wrenable_reg_22 <= 'X';
        wrenable_reg_23 <= 'X';
        wrenable_reg_24 <= 'X';
        wrenable_reg_25 <= 'X';
        wrenable_reg_26 <= 'X';
        wrenable_reg_27 <= 'X';
        wrenable_reg_28 <= 'X';
        wrenable_reg_29 <= 'X';
        wrenable_reg_3 <= 'X';
        wrenable_reg_30 <= 'X';
        wrenable_reg_31 <= 'X';
        wrenable_reg_32 <= 'X';
        wrenable_reg_33 <= 'X';
        wrenable_reg_34 <= 'X';
        wrenable_reg_35 <= 'X';
        wrenable_reg_36 <= 'X';
        wrenable_reg_37 <= 'X';
        wrenable_reg_38 <= 'X';
        wrenable_reg_39 <= 'X';
        wrenable_reg_4 <= 'X';
        wrenable_reg_40 <= 'X';
        wrenable_reg_41 <= 'X';
        wrenable_reg_42 <= 'X';
        wrenable_reg_43 <= 'X';
        wrenable_reg_44 <= 'X';
        wrenable_reg_45 <= 'X';
        wrenable_reg_46 <= 'X';
        wrenable_reg_47 <= 'X';
        wrenable_reg_5 <= 'X';
        wrenable_reg_6 <= 'X';
        wrenable_reg_7 <= 'X';
        wrenable_reg_8 <= 'X';
        wrenable_reg_9 <= 'X';
    end case;
  end process;

end controller_acc_0_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2022 Politecnico di Milano
-- Author(s): Marco Lattuada <marco.lattuada@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity flipflop_AR is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic;
  -- OUT
  out1 : out std_logic

);
end flipflop_AR;

architecture flipflop_AR_arch of flipflop_AR is
  
  signal reg_out1 : std_logic := '0';
  begin
    process(clock,reset)
    begin
      if(reset = '0') then
        reg_out1 <= '0';
      elsif(clock'event and clock = '1') then
        reg_out1 <= in1;
      end if;
    end process;
    out1 <= reg_out1;

end flipflop_AR_arch;

-- Top component for acc_0
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity acc_0b is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  param : in std_logic_vector(31 downto 0) ;
  result : in std_logic_vector(31 downto 0) ;
  M_Rdata_ram : in std_logic_vector(31 downto 0) ;
  M_DataRdy : in std_logic;
  Min_oe_ram : in std_logic;
  Min_we_ram : in std_logic;
  Min_addr_ram : in std_logic_vector(31 downto 0) ;
  Min_Wdata_ram : in std_logic_vector(31 downto 0) ;
  Min_data_ram_size : in std_logic_vector(5 downto 0) ;
  -- OUT
  done_port : out std_logic;
  Mout_oe_ram : out std_logic;
  Mout_we_ram : out std_logic;
  Mout_addr_ram : out std_logic_vector(31 downto 0) ;
  Mout_Wdata_ram : out std_logic_vector(31 downto 0) ;
  Mout_data_ram_size : out std_logic_vector(5 downto 0) 

);
end acc_0b;

architecture acc_0_archb of acc_0b is
  -- Component and signal declarations
  
  component datapath_acc_0
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in_port_param : in std_logic_vector(31 downto 0) ;
    in_port_result : in std_logic_vector(31 downto 0) ;
    M_Rdata_ram : in std_logic_vector(31 downto 0) ;
    M_DataRdy : in std_logic;
    Min_oe_ram : in std_logic;
    Min_we_ram : in std_logic;
    Min_addr_ram : in std_logic_vector(31 downto 0) ;
    Min_Wdata_ram : in std_logic_vector(31 downto 0) ;
    Min_data_ram_size : in std_logic_vector(5 downto 0) ;
    selector_IN_UNBOUNDED_acc_0_31017_31056 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31057 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31059 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31060 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31061 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31063 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31065 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31066 : in std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31068 : in std_logic;
    fuselector_MEMORY_CTRL_D21_251_i0_LOAD : in std_logic;
    fuselector_MEMORY_CTRL_D21_251_i0_STORE : in std_logic;
    selector_MUX_550_reg_13_0_0_0 : in std_logic;
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : in std_logic;
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : in std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : in std_logic;
    wrenable_reg_0 : in std_logic;
    wrenable_reg_1 : in std_logic;
    wrenable_reg_10 : in std_logic;
    wrenable_reg_11 : in std_logic;
    wrenable_reg_12 : in std_logic;
    wrenable_reg_13 : in std_logic;
    wrenable_reg_14 : in std_logic;
    wrenable_reg_15 : in std_logic;
    wrenable_reg_16 : in std_logic;
    wrenable_reg_17 : in std_logic;
    wrenable_reg_18 : in std_logic;
    wrenable_reg_19 : in std_logic;
    wrenable_reg_2 : in std_logic;
    wrenable_reg_20 : in std_logic;
    wrenable_reg_21 : in std_logic;
    wrenable_reg_22 : in std_logic;
    wrenable_reg_23 : in std_logic;
    wrenable_reg_24 : in std_logic;
    wrenable_reg_25 : in std_logic;
    wrenable_reg_26 : in std_logic;
    wrenable_reg_27 : in std_logic;
    wrenable_reg_28 : in std_logic;
    wrenable_reg_29 : in std_logic;
    wrenable_reg_3 : in std_logic;
    wrenable_reg_30 : in std_logic;
    wrenable_reg_31 : in std_logic;
    wrenable_reg_32 : in std_logic;
    wrenable_reg_33 : in std_logic;
    wrenable_reg_34 : in std_logic;
    wrenable_reg_35 : in std_logic;
    wrenable_reg_36 : in std_logic;
    wrenable_reg_37 : in std_logic;
    wrenable_reg_38 : in std_logic;
    wrenable_reg_39 : in std_logic;
    wrenable_reg_4 : in std_logic;
    wrenable_reg_40 : in std_logic;
    wrenable_reg_41 : in std_logic;
    wrenable_reg_42 : in std_logic;
    wrenable_reg_43 : in std_logic;
    wrenable_reg_44 : in std_logic;
    wrenable_reg_45 : in std_logic;
    wrenable_reg_46 : in std_logic;
    wrenable_reg_47 : in std_logic;
    wrenable_reg_5 : in std_logic;
    wrenable_reg_6 : in std_logic;
    wrenable_reg_7 : in std_logic;
    wrenable_reg_8 : in std_logic;
    wrenable_reg_9 : in std_logic;
    -- OUT
    Mout_oe_ram : out std_logic;
    Mout_we_ram : out std_logic;
    Mout_addr_ram : out std_logic_vector(31 downto 0) ;
    Mout_Wdata_ram : out std_logic_vector(31 downto 0) ;
    Mout_data_ram_size : out std_logic_vector(5 downto 0) ;
    OUT_MULTIIF_acc_0_31017_37300 : out std_logic_vector(0 downto 0);
    OUT_UNBOUNDED_acc_0_31017_31056 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31057 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31059 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31060 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31061 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31063 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31065 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31066 : out std_logic;
    OUT_UNBOUNDED_acc_0_31017_31068 : out std_logic
  
  );
  end component;
  
  component controller_acc_0
  port (
    -- IN
    OUT_MULTIIF_acc_0_31017_37300 : in std_logic_vector(0 downto 0);
    OUT_UNBOUNDED_acc_0_31017_31056 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31057 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31059 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31060 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31061 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31063 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31065 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31066 : in std_logic;
    OUT_UNBOUNDED_acc_0_31017_31068 : in std_logic;
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    -- OUT
    done_port : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31056 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31057 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31059 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31060 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31061 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31063 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31065 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31066 : out std_logic;
    selector_IN_UNBOUNDED_acc_0_31017_31068 : out std_logic;
    fuselector_MEMORY_CTRL_D21_251_i0_LOAD : out std_logic;
    fuselector_MEMORY_CTRL_D21_251_i0_STORE : out std_logic;
    selector_MUX_550_reg_13_0_0_0 : out std_logic;
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : out std_logic;
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : out std_logic;
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : out std_logic;
    wrenable_reg_0 : out std_logic;
    wrenable_reg_1 : out std_logic;
    wrenable_reg_10 : out std_logic;
    wrenable_reg_11 : out std_logic;
    wrenable_reg_12 : out std_logic;
    wrenable_reg_13 : out std_logic;
    wrenable_reg_14 : out std_logic;
    wrenable_reg_15 : out std_logic;
    wrenable_reg_16 : out std_logic;
    wrenable_reg_17 : out std_logic;
    wrenable_reg_18 : out std_logic;
    wrenable_reg_19 : out std_logic;
    wrenable_reg_2 : out std_logic;
    wrenable_reg_20 : out std_logic;
    wrenable_reg_21 : out std_logic;
    wrenable_reg_22 : out std_logic;
    wrenable_reg_23 : out std_logic;
    wrenable_reg_24 : out std_logic;
    wrenable_reg_25 : out std_logic;
    wrenable_reg_26 : out std_logic;
    wrenable_reg_27 : out std_logic;
    wrenable_reg_28 : out std_logic;
    wrenable_reg_29 : out std_logic;
    wrenable_reg_3 : out std_logic;
    wrenable_reg_30 : out std_logic;
    wrenable_reg_31 : out std_logic;
    wrenable_reg_32 : out std_logic;
    wrenable_reg_33 : out std_logic;
    wrenable_reg_34 : out std_logic;
    wrenable_reg_35 : out std_logic;
    wrenable_reg_36 : out std_logic;
    wrenable_reg_37 : out std_logic;
    wrenable_reg_38 : out std_logic;
    wrenable_reg_39 : out std_logic;
    wrenable_reg_4 : out std_logic;
    wrenable_reg_40 : out std_logic;
    wrenable_reg_41 : out std_logic;
    wrenable_reg_42 : out std_logic;
    wrenable_reg_43 : out std_logic;
    wrenable_reg_44 : out std_logic;
    wrenable_reg_45 : out std_logic;
    wrenable_reg_46 : out std_logic;
    wrenable_reg_47 : out std_logic;
    wrenable_reg_5 : out std_logic;
    wrenable_reg_6 : out std_logic;
    wrenable_reg_7 : out std_logic;
    wrenable_reg_8 : out std_logic;
    wrenable_reg_9 : out std_logic
  
  );
  end component;
  
  component flipflop_AR
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  signal OUT_MULTIIF_acc_0_31017_37300 : std_logic_vector(0 downto 0);
  signal OUT_UNBOUNDED_acc_0_31017_31056 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31057 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31059 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31060 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31061 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31063 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31065 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31066 : std_logic;
  signal OUT_UNBOUNDED_acc_0_31017_31068 : std_logic;
  signal done_delayed_REG_signal_in : std_logic;
  signal done_delayed_REG_signal_out : std_logic;
  signal fuselector_MEMORY_CTRL_D21_251_i0_LOAD : std_logic;
  signal fuselector_MEMORY_CTRL_D21_251_i0_STORE : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31056 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31057 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31059 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31060 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31061 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31063 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31065 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31066 : std_logic;
  signal selector_IN_UNBOUNDED_acc_0_31017_31068 : std_logic;
  signal selector_MUX_550_reg_13_0_0_0 : std_logic;
  signal selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 : std_logic;
  signal selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 : std_logic;
  signal selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 : std_logic;
  signal wrenable_reg_0 : std_logic;
  signal wrenable_reg_1 : std_logic;
  signal wrenable_reg_10 : std_logic;
  signal wrenable_reg_11 : std_logic;
  signal wrenable_reg_12 : std_logic;
  signal wrenable_reg_13 : std_logic;
  signal wrenable_reg_14 : std_logic;
  signal wrenable_reg_15 : std_logic;
  signal wrenable_reg_16 : std_logic;
  signal wrenable_reg_17 : std_logic;
  signal wrenable_reg_18 : std_logic;
  signal wrenable_reg_19 : std_logic;
  signal wrenable_reg_2 : std_logic;
  signal wrenable_reg_20 : std_logic;
  signal wrenable_reg_21 : std_logic;
  signal wrenable_reg_22 : std_logic;
  signal wrenable_reg_23 : std_logic;
  signal wrenable_reg_24 : std_logic;
  signal wrenable_reg_25 : std_logic;
  signal wrenable_reg_26 : std_logic;
  signal wrenable_reg_27 : std_logic;
  signal wrenable_reg_28 : std_logic;
  signal wrenable_reg_29 : std_logic;
  signal wrenable_reg_3 : std_logic;
  signal wrenable_reg_30 : std_logic;
  signal wrenable_reg_31 : std_logic;
  signal wrenable_reg_32 : std_logic;
  signal wrenable_reg_33 : std_logic;
  signal wrenable_reg_34 : std_logic;
  signal wrenable_reg_35 : std_logic;
  signal wrenable_reg_36 : std_logic;
  signal wrenable_reg_37 : std_logic;
  signal wrenable_reg_38 : std_logic;
  signal wrenable_reg_39 : std_logic;
  signal wrenable_reg_4 : std_logic;
  signal wrenable_reg_40 : std_logic;
  signal wrenable_reg_41 : std_logic;
  signal wrenable_reg_42 : std_logic;
  signal wrenable_reg_43 : std_logic;
  signal wrenable_reg_44 : std_logic;
  signal wrenable_reg_45 : std_logic;
  signal wrenable_reg_46 : std_logic;
  signal wrenable_reg_47 : std_logic;
  signal wrenable_reg_5 : std_logic;
  signal wrenable_reg_6 : std_logic;
  signal wrenable_reg_7 : std_logic;
  signal wrenable_reg_8 : std_logic;
  signal wrenable_reg_9 : std_logic;
begin
  Controller_i : controller_acc_0 port map (done_port => done_delayed_REG_signal_in,
    selector_IN_UNBOUNDED_acc_0_31017_31056 => selector_IN_UNBOUNDED_acc_0_31017_31056,
    selector_IN_UNBOUNDED_acc_0_31017_31057 => selector_IN_UNBOUNDED_acc_0_31017_31057,
    selector_IN_UNBOUNDED_acc_0_31017_31059 => selector_IN_UNBOUNDED_acc_0_31017_31059,
    selector_IN_UNBOUNDED_acc_0_31017_31060 => selector_IN_UNBOUNDED_acc_0_31017_31060,
    selector_IN_UNBOUNDED_acc_0_31017_31061 => selector_IN_UNBOUNDED_acc_0_31017_31061,
    selector_IN_UNBOUNDED_acc_0_31017_31063 => selector_IN_UNBOUNDED_acc_0_31017_31063,
    selector_IN_UNBOUNDED_acc_0_31017_31065 => selector_IN_UNBOUNDED_acc_0_31017_31065,
    selector_IN_UNBOUNDED_acc_0_31017_31066 => selector_IN_UNBOUNDED_acc_0_31017_31066,
    selector_IN_UNBOUNDED_acc_0_31017_31068 => selector_IN_UNBOUNDED_acc_0_31017_31068,
    fuselector_MEMORY_CTRL_D21_251_i0_LOAD => fuselector_MEMORY_CTRL_D21_251_i0_LOAD,
    fuselector_MEMORY_CTRL_D21_251_i0_STORE => fuselector_MEMORY_CTRL_D21_251_i0_STORE,
    selector_MUX_550_reg_13_0_0_0 => selector_MUX_550_reg_13_0_0_0,
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0,
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0,
    wrenable_reg_0 => wrenable_reg_0,
    wrenable_reg_1 => wrenable_reg_1,
    wrenable_reg_10 => wrenable_reg_10,
    wrenable_reg_11 => wrenable_reg_11,
    wrenable_reg_12 => wrenable_reg_12,
    wrenable_reg_13 => wrenable_reg_13,
    wrenable_reg_14 => wrenable_reg_14,
    wrenable_reg_15 => wrenable_reg_15,
    wrenable_reg_16 => wrenable_reg_16,
    wrenable_reg_17 => wrenable_reg_17,
    wrenable_reg_18 => wrenable_reg_18,
    wrenable_reg_19 => wrenable_reg_19,
    wrenable_reg_2 => wrenable_reg_2,
    wrenable_reg_20 => wrenable_reg_20,
    wrenable_reg_21 => wrenable_reg_21,
    wrenable_reg_22 => wrenable_reg_22,
    wrenable_reg_23 => wrenable_reg_23,
    wrenable_reg_24 => wrenable_reg_24,
    wrenable_reg_25 => wrenable_reg_25,
    wrenable_reg_26 => wrenable_reg_26,
    wrenable_reg_27 => wrenable_reg_27,
    wrenable_reg_28 => wrenable_reg_28,
    wrenable_reg_29 => wrenable_reg_29,
    wrenable_reg_3 => wrenable_reg_3,
    wrenable_reg_30 => wrenable_reg_30,
    wrenable_reg_31 => wrenable_reg_31,
    wrenable_reg_32 => wrenable_reg_32,
    wrenable_reg_33 => wrenable_reg_33,
    wrenable_reg_34 => wrenable_reg_34,
    wrenable_reg_35 => wrenable_reg_35,
    wrenable_reg_36 => wrenable_reg_36,
    wrenable_reg_37 => wrenable_reg_37,
    wrenable_reg_38 => wrenable_reg_38,
    wrenable_reg_39 => wrenable_reg_39,
    wrenable_reg_4 => wrenable_reg_4,
    wrenable_reg_40 => wrenable_reg_40,
    wrenable_reg_41 => wrenable_reg_41,
    wrenable_reg_42 => wrenable_reg_42,
    wrenable_reg_43 => wrenable_reg_43,
    wrenable_reg_44 => wrenable_reg_44,
    wrenable_reg_45 => wrenable_reg_45,
    wrenable_reg_46 => wrenable_reg_46,
    wrenable_reg_47 => wrenable_reg_47,
    wrenable_reg_5 => wrenable_reg_5,
    wrenable_reg_6 => wrenable_reg_6,
    wrenable_reg_7 => wrenable_reg_7,
    wrenable_reg_8 => wrenable_reg_8,
    wrenable_reg_9 => wrenable_reg_9,
    OUT_MULTIIF_acc_0_31017_37300 => OUT_MULTIIF_acc_0_31017_37300,
    OUT_UNBOUNDED_acc_0_31017_31056 => OUT_UNBOUNDED_acc_0_31017_31056,
    OUT_UNBOUNDED_acc_0_31017_31057 => OUT_UNBOUNDED_acc_0_31017_31057,
    OUT_UNBOUNDED_acc_0_31017_31059 => OUT_UNBOUNDED_acc_0_31017_31059,
    OUT_UNBOUNDED_acc_0_31017_31060 => OUT_UNBOUNDED_acc_0_31017_31060,
    OUT_UNBOUNDED_acc_0_31017_31061 => OUT_UNBOUNDED_acc_0_31017_31061,
    OUT_UNBOUNDED_acc_0_31017_31063 => OUT_UNBOUNDED_acc_0_31017_31063,
    OUT_UNBOUNDED_acc_0_31017_31065 => OUT_UNBOUNDED_acc_0_31017_31065,
    OUT_UNBOUNDED_acc_0_31017_31066 => OUT_UNBOUNDED_acc_0_31017_31066,
    OUT_UNBOUNDED_acc_0_31017_31068 => OUT_UNBOUNDED_acc_0_31017_31068,
    clock => clock,
    reset => reset,
    start_port => start_port);
  Datapath_i : datapath_acc_0 port map (Mout_oe_ram => Mout_oe_ram,
    Mout_we_ram => Mout_we_ram,
    Mout_addr_ram => Mout_addr_ram,
    Mout_Wdata_ram => Mout_Wdata_ram,
    Mout_data_ram_size => Mout_data_ram_size,
    OUT_MULTIIF_acc_0_31017_37300 => OUT_MULTIIF_acc_0_31017_37300,
    OUT_UNBOUNDED_acc_0_31017_31056 => OUT_UNBOUNDED_acc_0_31017_31056,
    OUT_UNBOUNDED_acc_0_31017_31057 => OUT_UNBOUNDED_acc_0_31017_31057,
    OUT_UNBOUNDED_acc_0_31017_31059 => OUT_UNBOUNDED_acc_0_31017_31059,
    OUT_UNBOUNDED_acc_0_31017_31060 => OUT_UNBOUNDED_acc_0_31017_31060,
    OUT_UNBOUNDED_acc_0_31017_31061 => OUT_UNBOUNDED_acc_0_31017_31061,
    OUT_UNBOUNDED_acc_0_31017_31063 => OUT_UNBOUNDED_acc_0_31017_31063,
    OUT_UNBOUNDED_acc_0_31017_31065 => OUT_UNBOUNDED_acc_0_31017_31065,
    OUT_UNBOUNDED_acc_0_31017_31066 => OUT_UNBOUNDED_acc_0_31017_31066,
    OUT_UNBOUNDED_acc_0_31017_31068 => OUT_UNBOUNDED_acc_0_31017_31068,
    clock => clock,
    reset => reset,
    in_port_param => param,
    in_port_result => result,
    M_Rdata_ram => M_Rdata_ram,
    M_DataRdy => M_DataRdy,
    Min_oe_ram => Min_oe_ram,
    Min_we_ram => Min_we_ram,
    Min_addr_ram => Min_addr_ram,
    Min_Wdata_ram => Min_Wdata_ram,
    Min_data_ram_size => Min_data_ram_size,
    selector_IN_UNBOUNDED_acc_0_31017_31056 => selector_IN_UNBOUNDED_acc_0_31017_31056,
    selector_IN_UNBOUNDED_acc_0_31017_31057 => selector_IN_UNBOUNDED_acc_0_31017_31057,
    selector_IN_UNBOUNDED_acc_0_31017_31059 => selector_IN_UNBOUNDED_acc_0_31017_31059,
    selector_IN_UNBOUNDED_acc_0_31017_31060 => selector_IN_UNBOUNDED_acc_0_31017_31060,
    selector_IN_UNBOUNDED_acc_0_31017_31061 => selector_IN_UNBOUNDED_acc_0_31017_31061,
    selector_IN_UNBOUNDED_acc_0_31017_31063 => selector_IN_UNBOUNDED_acc_0_31017_31063,
    selector_IN_UNBOUNDED_acc_0_31017_31065 => selector_IN_UNBOUNDED_acc_0_31017_31065,
    selector_IN_UNBOUNDED_acc_0_31017_31066 => selector_IN_UNBOUNDED_acc_0_31017_31066,
    selector_IN_UNBOUNDED_acc_0_31017_31068 => selector_IN_UNBOUNDED_acc_0_31017_31068,
    fuselector_MEMORY_CTRL_D21_251_i0_LOAD => fuselector_MEMORY_CTRL_D21_251_i0_LOAD,
    fuselector_MEMORY_CTRL_D21_251_i0_STORE => fuselector_MEMORY_CTRL_D21_251_i0_STORE,
    selector_MUX_550_reg_13_0_0_0 => selector_MUX_550_reg_13_0_0_0,
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0 => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_0,
    selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1 => selector_MUX_5_MEMORY_CTRL_D21_251_i0_0_0_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_0,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_2,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_3,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_0_4,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_0,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_1,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_1_2,
    selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0 => selector_MUX_6_MEMORY_CTRL_D21_251_i0_1_2_0,
    wrenable_reg_0 => wrenable_reg_0,
    wrenable_reg_1 => wrenable_reg_1,
    wrenable_reg_10 => wrenable_reg_10,
    wrenable_reg_11 => wrenable_reg_11,
    wrenable_reg_12 => wrenable_reg_12,
    wrenable_reg_13 => wrenable_reg_13,
    wrenable_reg_14 => wrenable_reg_14,
    wrenable_reg_15 => wrenable_reg_15,
    wrenable_reg_16 => wrenable_reg_16,
    wrenable_reg_17 => wrenable_reg_17,
    wrenable_reg_18 => wrenable_reg_18,
    wrenable_reg_19 => wrenable_reg_19,
    wrenable_reg_2 => wrenable_reg_2,
    wrenable_reg_20 => wrenable_reg_20,
    wrenable_reg_21 => wrenable_reg_21,
    wrenable_reg_22 => wrenable_reg_22,
    wrenable_reg_23 => wrenable_reg_23,
    wrenable_reg_24 => wrenable_reg_24,
    wrenable_reg_25 => wrenable_reg_25,
    wrenable_reg_26 => wrenable_reg_26,
    wrenable_reg_27 => wrenable_reg_27,
    wrenable_reg_28 => wrenable_reg_28,
    wrenable_reg_29 => wrenable_reg_29,
    wrenable_reg_3 => wrenable_reg_3,
    wrenable_reg_30 => wrenable_reg_30,
    wrenable_reg_31 => wrenable_reg_31,
    wrenable_reg_32 => wrenable_reg_32,
    wrenable_reg_33 => wrenable_reg_33,
    wrenable_reg_34 => wrenable_reg_34,
    wrenable_reg_35 => wrenable_reg_35,
    wrenable_reg_36 => wrenable_reg_36,
    wrenable_reg_37 => wrenable_reg_37,
    wrenable_reg_38 => wrenable_reg_38,
    wrenable_reg_39 => wrenable_reg_39,
    wrenable_reg_4 => wrenable_reg_4,
    wrenable_reg_40 => wrenable_reg_40,
    wrenable_reg_41 => wrenable_reg_41,
    wrenable_reg_42 => wrenable_reg_42,
    wrenable_reg_43 => wrenable_reg_43,
    wrenable_reg_44 => wrenable_reg_44,
    wrenable_reg_45 => wrenable_reg_45,
    wrenable_reg_46 => wrenable_reg_46,
    wrenable_reg_47 => wrenable_reg_47,
    wrenable_reg_5 => wrenable_reg_5,
    wrenable_reg_6 => wrenable_reg_6,
    wrenable_reg_7 => wrenable_reg_7,
    wrenable_reg_8 => wrenable_reg_8,
    wrenable_reg_9 => wrenable_reg_9);
  done_delayed_REG : flipflop_AR generic map(BITSIZE_in1=>1,
    BITSIZE_out1=>1) port map (out1 => done_delayed_REG_signal_out,
    clock => clock,
    reset => reset,
    in1 => done_delayed_REG_signal_in);
  -- io-signal post fix
  done_port <= done_delayed_REG_signal_out;

end acc_0_archb;

-- Minimal interface for function: acc_0
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity acc_0 is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  param : in std_logic_vector(31 downto 0) ;
  result : in std_logic_vector(31 downto 0) ;
  M_Rdata_ram : in std_logic_vector(31 downto 0) ;
  M_DataRdy : in std_logic;
  -- OUT
  done_port : out std_logic;
  Mout_oe_ram : out std_logic;
  Mout_we_ram : out std_logic;
  Mout_addr_ram : out std_logic_vector(31 downto 0) ;
  Mout_Wdata_ram : out std_logic_vector(31 downto 0) ;
  Mout_data_ram_size : out std_logic_vector(5 downto 0) 

);
end acc_0;

architecture acc_0_arch of acc_0 is
  -- Component and signal declarations
  
  component acc_0b
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    param : in std_logic_vector(31 downto 0) ;
    result : in std_logic_vector(31 downto 0) ;
    M_Rdata_ram : in std_logic_vector(31 downto 0) ;
    M_DataRdy : in std_logic;
    Min_oe_ram : in std_logic;
    Min_we_ram : in std_logic;
    Min_addr_ram : in std_logic_vector(31 downto 0) ;
    Min_Wdata_ram : in std_logic_vector(31 downto 0) ;
    Min_data_ram_size : in std_logic_vector(5 downto 0) ;
    -- OUT
    done_port : out std_logic;
    Mout_oe_ram : out std_logic;
    Mout_we_ram : out std_logic;
    Mout_addr_ram : out std_logic_vector(31 downto 0) ;
    Mout_Wdata_ram : out std_logic_vector(31 downto 0) ;
    Mout_data_ram_size : out std_logic_vector(5 downto 0) 
  
  );
  end component;
begin
  \_acc_0_i0\ : acc_0b port map (done_port => done_port,
    Mout_oe_ram => Mout_oe_ram,
    Mout_we_ram => Mout_we_ram,
    Mout_addr_ram => Mout_addr_ram,
    Mout_Wdata_ram => Mout_Wdata_ram,
    Mout_data_ram_size => Mout_data_ram_size,
    clock => clock,
    reset => reset,
    start_port => start_port,
    param => param,
    result => result,
    M_Rdata_ram => M_Rdata_ram,
    M_DataRdy => M_DataRdy,
    Min_oe_ram => '0',
    Min_we_ram => '0',
    Min_addr_ram => "00000000000000000000000000000000",
    Min_Wdata_ram => "00000000000000000000000000000000",
    Min_data_ram_size => "000000");

end acc_0_arch;


